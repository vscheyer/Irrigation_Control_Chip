magic
tech sky130A
timestamp 1619709734
<< nwell >>
rect 18710 1340 20015 1545
<< nmos >>
rect 19495 1205 19995 1255
rect 18845 1095 18860 1195
rect 18910 1095 18925 1195
rect 19060 1095 19075 1195
rect 19210 1095 19225 1195
<< pmos >>
rect 18845 1395 18860 1495
rect 18910 1395 18925 1495
rect 19060 1395 19075 1495
rect 19210 1395 19225 1495
rect 19495 1420 19995 1470
<< ndiff >>
rect 19495 1290 19995 1305
rect 19495 1270 19510 1290
rect 19980 1270 19995 1290
rect 19495 1255 19995 1270
rect 18795 1185 18845 1195
rect 18795 1105 18810 1185
rect 18830 1105 18845 1185
rect 18795 1095 18845 1105
rect 18860 1185 18910 1195
rect 18860 1105 18875 1185
rect 18895 1105 18910 1185
rect 18860 1095 18910 1105
rect 18925 1185 18975 1195
rect 18925 1105 18940 1185
rect 18960 1105 18975 1185
rect 18925 1095 18975 1105
rect 19010 1185 19060 1195
rect 19010 1105 19025 1185
rect 19045 1105 19060 1185
rect 19010 1095 19060 1105
rect 19075 1185 19125 1195
rect 19075 1105 19090 1185
rect 19110 1105 19125 1185
rect 19075 1095 19125 1105
rect 19160 1185 19210 1195
rect 19160 1105 19175 1185
rect 19195 1105 19210 1185
rect 19160 1095 19210 1105
rect 19225 1185 19275 1195
rect 19225 1105 19240 1185
rect 19260 1105 19275 1185
rect 19495 1190 19995 1205
rect 19495 1170 19510 1190
rect 19980 1170 19995 1190
rect 19495 1155 19995 1170
rect 19225 1095 19275 1105
<< pdiff >>
rect 19495 1505 19995 1520
rect 18795 1485 18845 1495
rect 18795 1405 18810 1485
rect 18830 1405 18845 1485
rect 18795 1395 18845 1405
rect 18860 1485 18910 1495
rect 18860 1405 18875 1485
rect 18895 1405 18910 1485
rect 18860 1395 18910 1405
rect 18925 1485 18975 1495
rect 18925 1405 18940 1485
rect 18960 1405 18975 1485
rect 18925 1395 18975 1405
rect 19010 1485 19060 1495
rect 19010 1405 19025 1485
rect 19045 1405 19060 1485
rect 19010 1395 19060 1405
rect 19075 1485 19125 1495
rect 19075 1405 19090 1485
rect 19110 1405 19125 1485
rect 19075 1395 19125 1405
rect 19160 1485 19210 1495
rect 19160 1405 19175 1485
rect 19195 1405 19210 1485
rect 19160 1395 19210 1405
rect 19225 1485 19275 1495
rect 19225 1405 19240 1485
rect 19260 1405 19275 1485
rect 19495 1485 19510 1505
rect 19980 1485 19995 1505
rect 19495 1470 19995 1485
rect 19225 1395 19275 1405
rect 19495 1405 19995 1420
rect 19495 1385 19510 1405
rect 19980 1385 19995 1405
rect 19495 1370 19995 1385
<< ndiffc >>
rect 19510 1270 19980 1290
rect 18810 1105 18830 1185
rect 18875 1105 18895 1185
rect 18940 1105 18960 1185
rect 19025 1105 19045 1185
rect 19090 1105 19110 1185
rect 19175 1105 19195 1185
rect 19240 1105 19260 1185
rect 19510 1170 19980 1190
<< pdiffc >>
rect 18810 1405 18830 1485
rect 18875 1405 18895 1485
rect 18940 1405 18960 1485
rect 19025 1405 19045 1485
rect 19090 1405 19110 1485
rect 19175 1405 19195 1485
rect 19240 1405 19260 1485
rect 19510 1485 19980 1505
rect 19510 1385 19980 1405
<< psubdiff >>
rect 20065 1535 20115 1545
rect 20065 1455 20080 1535
rect 20100 1455 20115 1535
rect 20065 1445 20115 1455
rect 18745 1185 18795 1195
rect 18745 1105 18760 1185
rect 18780 1105 18795 1185
rect 18745 1095 18795 1105
<< nsubdiff >>
rect 18745 1485 18795 1495
rect 18745 1405 18760 1485
rect 18780 1405 18795 1485
rect 18745 1395 18795 1405
<< psubdiffcont >>
rect 20080 1455 20100 1535
rect 18760 1105 18780 1185
<< nsubdiffcont >>
rect 18760 1405 18780 1485
<< poly >>
rect 18820 1540 18860 1550
rect 18820 1520 18830 1540
rect 18850 1520 18860 1540
rect 18820 1510 18860 1520
rect 19060 1540 19100 1550
rect 19060 1520 19070 1540
rect 19090 1520 19100 1540
rect 19060 1510 19100 1520
rect 18845 1495 18860 1510
rect 18910 1495 18925 1510
rect 19060 1495 19075 1510
rect 19210 1495 19225 1510
rect 19470 1420 19495 1470
rect 19995 1420 20010 1470
rect 18845 1385 18860 1395
rect 18910 1385 18925 1395
rect 18845 1370 18925 1385
rect 18845 1220 18860 1370
rect 18910 1220 18925 1370
rect 19060 1315 19075 1395
rect 19035 1305 19075 1315
rect 19035 1285 19045 1305
rect 19065 1290 19075 1305
rect 19210 1290 19225 1395
rect 19470 1355 19485 1420
rect 19445 1345 19485 1355
rect 19445 1325 19455 1345
rect 19475 1325 19485 1345
rect 19445 1315 19485 1325
rect 19065 1285 19225 1290
rect 19035 1275 19225 1285
rect 18845 1205 18925 1220
rect 18845 1195 18860 1205
rect 18910 1195 18925 1205
rect 19060 1195 19075 1275
rect 19210 1195 19225 1275
rect 19470 1255 19485 1315
rect 19470 1205 19495 1255
rect 19995 1205 20010 1255
rect 18845 1080 18860 1095
rect 18910 1080 18925 1095
rect 19060 1080 19075 1095
rect 19210 1080 19225 1095
<< polycont >>
rect 18830 1520 18850 1540
rect 19070 1520 19090 1540
rect 19045 1285 19065 1305
rect 19455 1325 19475 1345
<< xpolycontact >>
rect 18690 3570 18725 3790
rect 18690 1600 18725 1820
rect 18850 3570 18885 3790
rect 18850 1600 18885 1820
rect 19010 3570 19045 3790
rect 19010 1600 19045 1820
rect 19170 3570 19205 3790
rect 19170 1600 19205 1820
rect 19330 3570 19365 3790
rect 19330 1600 19365 1820
rect 19490 3570 19525 3790
rect 19490 1600 19525 1820
rect 19650 3570 19685 3790
rect 19650 1600 19685 1820
rect 19810 3570 19845 3790
rect 19810 1600 19845 1820
rect 19970 3570 20005 3790
rect 19970 1600 20005 1820
rect 20130 3570 20165 3790
rect 20130 1600 20165 1820
<< xpolyres >>
rect 18690 1820 18725 3570
rect 18850 1820 18885 3570
rect 19010 1820 19045 3570
rect 19170 1820 19205 3570
rect 19330 1820 19365 3570
rect 19490 1820 19525 3570
rect 19650 1820 19685 3570
rect 19810 1820 19845 3570
rect 19970 1820 20005 3570
rect 20130 1820 20165 3570
<< locali >>
rect 18725 3570 18850 3790
rect 19045 3570 19170 3790
rect 19365 3570 19490 3790
rect 19685 3570 19810 3790
rect 20005 3570 20130 3790
rect 18885 1600 19010 1820
rect 19205 1600 19330 1820
rect 19525 1600 19650 1820
rect 19845 1600 19970 1820
rect 18690 1550 18725 1600
rect 20130 1580 20165 1600
rect 19080 1560 20165 1580
rect 19080 1550 19100 1560
rect 18690 1540 18860 1550
rect 18690 1530 18830 1540
rect 18820 1520 18830 1530
rect 18850 1520 18860 1540
rect 19060 1540 19100 1550
rect 18820 1510 18860 1520
rect 18885 1510 19035 1530
rect 19060 1520 19070 1540
rect 19090 1520 19100 1540
rect 19060 1510 19100 1520
rect 20070 1535 20110 1540
rect 18885 1490 18905 1510
rect 19015 1490 19035 1510
rect 19500 1505 19990 1515
rect 18750 1485 18840 1490
rect 18750 1405 18760 1485
rect 18780 1405 18810 1485
rect 18830 1405 18840 1485
rect 18750 1400 18840 1405
rect 18865 1485 18905 1490
rect 18865 1405 18875 1485
rect 18895 1405 18905 1485
rect 18865 1400 18905 1405
rect 18930 1485 18970 1490
rect 18930 1405 18940 1485
rect 18960 1405 18970 1485
rect 18930 1400 18970 1405
rect 19015 1485 19055 1490
rect 19015 1405 19025 1485
rect 19045 1405 19055 1485
rect 19015 1400 19055 1405
rect 19080 1485 19120 1490
rect 19080 1405 19090 1485
rect 19110 1405 19120 1485
rect 19080 1400 19120 1405
rect 19165 1485 19205 1490
rect 19165 1405 19175 1485
rect 19195 1405 19205 1485
rect 19165 1400 19205 1405
rect 19230 1485 19270 1490
rect 19230 1405 19240 1485
rect 19260 1405 19270 1485
rect 19500 1485 19510 1505
rect 19980 1485 19990 1505
rect 19500 1475 19990 1485
rect 20070 1455 20080 1535
rect 20100 1455 20110 1535
rect 20070 1450 20110 1455
rect 19230 1400 19270 1405
rect 18930 1295 18950 1400
rect 19250 1335 19270 1400
rect 19500 1405 20165 1415
rect 19500 1385 19510 1405
rect 19980 1395 20165 1405
rect 19980 1385 19990 1395
rect 19500 1375 19990 1385
rect 19445 1345 19485 1355
rect 19445 1335 19455 1345
rect 19250 1325 19455 1335
rect 19475 1325 19485 1345
rect 19250 1315 19485 1325
rect 19035 1305 19075 1315
rect 19035 1295 19045 1305
rect 18690 1285 19045 1295
rect 19065 1285 19075 1305
rect 18690 1275 19075 1285
rect 18930 1190 18950 1275
rect 18970 1245 19020 1255
rect 18970 1220 18975 1245
rect 19015 1240 19020 1245
rect 19015 1220 19100 1240
rect 18970 1210 19020 1220
rect 19080 1190 19100 1220
rect 19250 1190 19270 1315
rect 19970 1300 19990 1375
rect 19500 1290 19990 1300
rect 19500 1270 19510 1290
rect 19980 1270 19990 1290
rect 19500 1260 19990 1270
rect 18750 1185 18840 1190
rect 18750 1105 18760 1185
rect 18780 1105 18810 1185
rect 18830 1105 18840 1185
rect 18750 1100 18840 1105
rect 18865 1185 18905 1190
rect 18865 1105 18875 1185
rect 18895 1105 18905 1185
rect 18865 1100 18905 1105
rect 18930 1185 18970 1190
rect 18930 1105 18940 1185
rect 18960 1105 18970 1185
rect 18930 1100 18970 1105
rect 19015 1185 19055 1190
rect 19015 1105 19025 1185
rect 19045 1105 19055 1185
rect 19015 1100 19055 1105
rect 19080 1185 19120 1190
rect 19080 1105 19090 1185
rect 19110 1105 19120 1185
rect 19080 1100 19120 1105
rect 19165 1185 19205 1190
rect 19165 1105 19175 1185
rect 19195 1105 19205 1185
rect 19165 1100 19205 1105
rect 19230 1185 19270 1190
rect 19230 1105 19240 1185
rect 19260 1105 19270 1185
rect 19500 1190 19990 1200
rect 19500 1170 19510 1190
rect 19980 1170 19990 1190
rect 19500 1160 19990 1170
rect 19230 1100 19270 1105
rect 18885 1080 18905 1100
rect 19015 1080 19035 1100
rect 18885 1060 19035 1080
<< viali >>
rect 18760 1405 18780 1485
rect 18810 1405 18830 1485
rect 19090 1405 19110 1485
rect 19175 1405 19195 1485
rect 19510 1485 19980 1505
rect 18975 1220 19015 1245
rect 18760 1105 18780 1185
rect 18810 1105 18830 1185
rect 19175 1105 19195 1185
rect 19510 1170 19980 1190
<< metal1 >>
rect 18800 1515 19205 1520
rect 18800 1505 19990 1515
rect 18800 1490 18840 1505
rect 18690 1485 18840 1490
rect 18690 1405 18760 1485
rect 18780 1405 18810 1485
rect 18830 1405 18840 1485
rect 18690 1400 18840 1405
rect 18750 1255 18840 1400
rect 19035 1485 19120 1490
rect 19035 1405 19090 1485
rect 19110 1405 19120 1485
rect 19035 1400 19120 1405
rect 19165 1485 19510 1505
rect 19980 1485 19990 1505
rect 19165 1405 19175 1485
rect 19195 1475 19990 1485
rect 19195 1405 19205 1475
rect 19165 1400 19205 1405
rect 18750 1245 19020 1255
rect 18750 1220 18975 1245
rect 19015 1220 19020 1245
rect 18750 1210 19020 1220
rect 18750 1205 19005 1210
rect 19035 1190 19055 1400
rect 20070 1200 20110 1540
rect 19500 1190 20110 1200
rect 18690 1185 19510 1190
rect 18690 1105 18760 1185
rect 18780 1105 18810 1185
rect 18830 1105 19175 1185
rect 19195 1170 19510 1185
rect 19980 1170 20110 1190
rect 19195 1160 20110 1170
rect 19195 1105 19205 1160
rect 18690 1100 19205 1105
<< labels >>
rlabel metal1 18690 1445 18690 1445 7 VP
rlabel metal1 18690 1145 18690 1145 7 VN
rlabel locali 18690 1540 18690 1540 7 crystal1
rlabel locali 18690 1285 18690 1285 7 crystal2
rlabel locali 20165 1405 20165 1405 3 clk
<< end >>
