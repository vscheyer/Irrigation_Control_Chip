magic
tech sky130A
timestamp 1620791811
<< locali >>
rect -15360 17715 -15280 17725
rect -15360 17695 -15350 17715
rect -15290 17695 -15280 17715
rect -15460 17610 -15380 17620
rect -15460 17590 -15450 17610
rect -15390 17590 -15380 17610
rect -15460 13700 -15380 17590
rect -15460 13680 -15450 13700
rect -15390 13680 -15380 13700
rect -15460 9855 -15380 13680
rect -15360 13805 -15280 17695
rect -15360 13785 -15350 13805
rect -15290 13785 -15280 13805
rect -15360 9960 -15280 13785
rect -15360 9940 -15350 9960
rect -15290 9940 -15280 9960
rect -15360 9930 -15280 9940
rect -15460 9835 -15450 9855
rect -15390 9835 -15380 9855
rect -15460 9825 -15380 9835
<< viali >>
rect -15350 17695 -15290 17715
rect -15450 17590 -15390 17610
rect -15450 13680 -15390 13700
rect -15350 13785 -15290 13805
rect -15350 9940 -15290 9960
rect -15450 9835 -15390 9855
<< metal1 >>
rect -6500 19260 -6370 19350
rect -6500 17855 -6460 19260
rect -4970 19020 -4690 19060
rect -15360 17715 -15280 17725
rect -15360 17695 -15350 17715
rect -15290 17695 -15280 17715
rect -15360 17685 -15280 17695
rect -4730 16865 -4690 19020
rect -4935 16825 -4690 16865
rect -15360 13805 -15280 13815
rect -15360 13785 -15350 13805
rect -15290 13785 -15280 13805
rect -15360 13775 -15280 13785
rect -15360 9960 -15280 9970
rect -15360 9940 -15350 9960
rect -15290 9940 -15280 9960
rect -15360 9930 -15280 9940
use anADC  anADC_0
timestamp 1620787225
transform 1 0 -5702 0 1 10017
box -10150 -2930 995 145
use anADC  anADC_1
timestamp 1620787225
transform 1 0 -5702 0 1 13860
box -10150 -2930 995 145
use anADC  anADC_2
timestamp 1620787225
transform 1 0 -5735 0 1 17771
box -10150 -2930 995 145
use clock  clock_0
timestamp 1619709734
transform 1 0 -25069 0 1 17860
box 18690 1060 20165 3790
use fsm  fsm_0
timestamp 1620791022
transform 1 0 -2704 0 1 6075
box 0 0 15012 16084
<< end >>
