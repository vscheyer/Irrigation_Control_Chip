magic
tech sky130A
timestamp 1620637795
<< nwell >>
rect -7865 80 -7485 115
rect -7865 -10 -7455 80
rect -4840 70 -4380 115
rect -7865 -45 -7485 -10
rect -4855 -45 -4770 70
rect -4435 65 -4380 70
rect -4525 -25 -4380 65
rect -4855 -55 -4700 -45
rect -4850 -60 -4700 -55
rect -4435 -60 -4380 -25
rect -4275 -75 -4235 -50
rect -7490 -110 -7315 -75
rect -1780 -210 -1630 115
rect -4410 -350 -4405 -210
rect -1795 -350 -1630 -210
rect -1780 -375 -1630 -350
rect 625 -1190 965 -985
<< nmos >>
rect -7740 -220 -7725 -120
rect -7590 -220 -7575 -120
rect 240 -1070 540 -1055
<< pmos >>
rect -7740 -15 -7725 85
rect -7590 -15 -7575 85
rect 645 -1070 945 -1055
<< ndiff >>
rect -7790 -135 -7740 -120
rect -7790 -205 -7775 -135
rect -7755 -205 -7740 -135
rect -7790 -220 -7740 -205
rect -7725 -135 -7675 -120
rect -7725 -205 -7710 -135
rect -7690 -205 -7675 -135
rect -7725 -220 -7675 -205
rect -7640 -135 -7590 -120
rect -7640 -205 -7625 -135
rect -7605 -205 -7590 -135
rect -7640 -220 -7590 -205
rect -7575 -135 -7525 -120
rect -7575 -205 -7560 -135
rect -7540 -205 -7525 -135
rect -7575 -220 -7525 -205
rect 240 -1020 540 -1005
rect 240 -1040 255 -1020
rect 525 -1040 540 -1020
rect 240 -1055 540 -1040
rect 240 -1085 540 -1070
rect 240 -1105 255 -1085
rect 525 -1105 540 -1085
rect 240 -1120 540 -1105
<< pdiff >>
rect -7790 70 -7740 85
rect -7790 0 -7775 70
rect -7755 0 -7740 70
rect -7790 -15 -7740 0
rect -7725 70 -7675 85
rect -7725 0 -7710 70
rect -7690 0 -7675 70
rect -7725 -15 -7675 0
rect -7640 70 -7590 85
rect -7640 0 -7625 70
rect -7605 0 -7590 70
rect -7640 -15 -7590 0
rect -7575 70 -7525 85
rect -7575 0 -7560 70
rect -7540 0 -7525 70
rect -7575 -15 -7525 0
rect 645 -1020 945 -1005
rect 645 -1040 660 -1020
rect 930 -1040 945 -1020
rect 645 -1055 945 -1040
rect 645 -1085 945 -1070
rect 645 -1105 660 -1085
rect 930 -1105 945 -1085
rect 645 -1120 945 -1105
<< ndiffc >>
rect -7775 -205 -7755 -135
rect -7710 -205 -7690 -135
rect -7625 -205 -7605 -135
rect -7560 -205 -7540 -135
rect -4660 -220 -4640 -150
rect 255 -1040 525 -1020
rect 255 -1105 525 -1085
<< pdiffc >>
rect -7775 0 -7755 70
rect -7710 0 -7690 70
rect -7625 0 -7605 70
rect -7560 0 -7540 70
rect 660 -1040 930 -1020
rect 660 -1105 930 -1085
<< psubdiff >>
rect -5330 -2315 -5180 -2300
rect -5330 -2335 -5315 -2315
rect -5195 -2335 -5180 -2315
rect -5330 -2350 -5180 -2335
<< nsubdiff >>
rect 645 -1135 945 -1120
rect 645 -1155 660 -1135
rect 930 -1155 945 -1135
rect 645 -1170 945 -1155
<< psubdiffcont >>
rect -5315 -2335 -5195 -2315
<< nsubdiffcont >>
rect 660 -1155 930 -1135
<< poly >>
rect -7740 85 -7725 100
rect -7590 85 -7575 145
rect -4545 75 -4530 145
rect -7740 -30 -7725 -15
rect -7740 -40 -7615 -30
rect -7740 -45 -7645 -40
rect -7655 -60 -7645 -45
rect -7625 -60 -7615 -40
rect -7655 -70 -7615 -60
rect -7740 -120 -7725 -105
rect -7590 -120 -7575 -15
rect -7740 -230 -7725 -220
rect -7590 -230 -7575 -220
rect -7740 -245 -7575 -230
rect 955 -830 995 -820
rect 955 -850 965 -830
rect 985 -850 995 -830
rect 955 -860 995 -850
rect 955 -1055 970 -860
rect 225 -1070 240 -1055
rect 540 -1070 645 -1055
rect 945 -1070 970 -1055
<< polycont >>
rect -7645 -60 -7625 -40
rect 965 -850 985 -830
<< xpolycontact >>
rect -4415 -1155 -4195 -1120
rect -2005 -1155 -1785 -1120
rect -4415 -1315 -4195 -1280
rect -2005 -1315 -1785 -1280
rect -4415 -1475 -4195 -1440
rect -2005 -1475 -1785 -1440
rect -4415 -1635 -4195 -1600
rect -2005 -1635 -1785 -1600
rect -4415 -1795 -4195 -1760
rect -2005 -1795 -1785 -1760
rect -4415 -1955 -4195 -1920
rect -2005 -1955 -1785 -1920
rect -4415 -2115 -4195 -2080
rect -2005 -2115 -1785 -2080
rect -4415 -2275 -4195 -2240
rect -2005 -2275 -1785 -2240
rect -10150 -2435 -9930 -2400
rect -5080 -2435 -4860 -2400
rect -4735 -2435 -4515 -2400
rect 775 -2435 995 -2400
rect -10150 -2600 -9930 -2565
rect -5080 -2600 -4860 -2565
rect -4735 -2600 -4515 -2565
rect 775 -2600 995 -2565
rect -10150 -2765 -9930 -2730
rect -5080 -2765 -4860 -2730
rect -4735 -2765 -4515 -2730
rect 775 -2765 995 -2730
rect -10150 -2930 -9930 -2895
rect -5080 -2930 -4860 -2895
rect -4735 -2930 -4515 -2895
rect 775 -2930 995 -2895
<< xpolyres >>
rect -4195 -1155 -2005 -1120
rect -4195 -1315 -2005 -1280
rect -4195 -1475 -2005 -1440
rect -4195 -1635 -2005 -1600
rect -4195 -1795 -2005 -1760
rect -4195 -1955 -2005 -1920
rect -4195 -2115 -2005 -2080
rect -4195 -2275 -2005 -2240
rect -9930 -2435 -5080 -2400
rect -4515 -2435 775 -2400
rect -9930 -2600 -5080 -2565
rect -4515 -2600 775 -2565
rect -9930 -2765 -5080 -2730
rect -4515 -2765 775 -2730
rect -9930 -2930 -5080 -2895
rect -4515 -2930 775 -2895
<< locali >>
rect -7840 -85 -7820 145
rect -7870 -105 -7820 -85
rect -7785 70 -7745 80
rect -7785 0 -7775 70
rect -7755 0 -7745 70
rect -7785 -135 -7745 0
rect -7785 -205 -7775 -135
rect -7755 -205 -7745 -135
rect -7785 -215 -7745 -205
rect -7720 70 -7680 80
rect -7720 0 -7710 70
rect -7690 0 -7680 70
rect -7720 -135 -7680 0
rect -7635 70 -7595 80
rect -7635 0 -7625 70
rect -7605 0 -7595 70
rect -7635 -10 -7595 0
rect -7570 70 -7530 80
rect -7570 0 -7560 70
rect -7540 0 -7530 70
rect -7570 -10 -7530 0
rect -4525 55 -4435 65
rect -7635 -30 -7615 -10
rect -4525 -15 -4515 55
rect -4495 -15 -4465 55
rect -4445 -15 -4435 55
rect -4525 -25 -4435 -15
rect -4425 -25 -4390 65
rect -1765 -10 -1745 145
rect -7655 -40 -7615 -30
rect -7655 -60 -7645 -40
rect -7625 -60 -7615 -40
rect -7655 -70 -7615 -60
rect -7720 -205 -7710 -135
rect -7690 -205 -7680 -135
rect -8190 -255 -8170 -225
rect -7785 -255 -7765 -215
rect -8190 -275 -7765 -255
rect -7720 -245 -7680 -205
rect -7635 -125 -7615 -70
rect -4425 -120 -4410 -100
rect -7635 -135 -7595 -125
rect -7635 -205 -7625 -135
rect -7605 -205 -7595 -135
rect -7635 -215 -7595 -205
rect -7570 -135 -7530 -125
rect -7570 -205 -7560 -135
rect -7540 -205 -7530 -135
rect -7570 -215 -7530 -205
rect -4420 -230 -4410 -140
rect -7720 -275 -7500 -245
rect -7580 -405 -7500 -275
rect -4735 -270 -4715 -240
rect -4670 -250 -4650 -240
rect -4735 -290 -4485 -270
rect -7580 -425 -7570 -405
rect -7510 -425 -7500 -405
rect -7580 -435 -7500 -425
rect -4905 -400 -4825 -390
rect -4905 -420 -4895 -400
rect -4835 -420 -4825 -400
rect -4905 -430 -4825 -420
rect -7560 -505 -7520 -495
rect -7560 -565 -7550 -505
rect -7530 -565 -7520 -505
rect -7560 -1070 -7520 -565
rect -4830 -860 -4525 -840
rect -4830 -900 -4695 -880
rect -7560 -1110 -7330 -1070
rect -7370 -1370 -7330 -1110
rect -4715 -1245 -4695 -900
rect -4715 -1255 -4565 -1245
rect -7475 -1380 -7325 -1370
rect -7475 -1620 -7465 -1380
rect -7335 -1620 -7325 -1380
rect -4715 -1495 -4705 -1255
rect -4575 -1495 -4565 -1255
rect -4715 -1505 -4565 -1495
rect -7475 -1630 -7325 -1620
rect -4545 -1650 -4525 -860
rect -4715 -1660 -4525 -1650
rect -4715 -1900 -4705 -1660
rect -4575 -1670 -4525 -1660
rect -4505 -1175 -4485 -290
rect -4465 -505 -4385 -495
rect -4465 -525 -4455 -505
rect -4395 -525 -4385 -505
rect -4465 -535 -4385 -525
rect -1750 -505 -1645 -495
rect -1750 -525 -1715 -505
rect -1655 -525 -1645 -505
rect -1750 -535 -1645 -525
rect -4465 -1120 -4445 -535
rect -1745 -860 -1670 -535
rect 955 -830 995 -820
rect 955 -850 965 -830
rect 985 -850 995 -830
rect 955 -860 995 -850
rect -4465 -1155 -4415 -1120
rect -4575 -1900 -4565 -1670
rect -4715 -1910 -4565 -1900
rect -4505 -2240 -4435 -1175
rect -4415 -1440 -4195 -1315
rect -4415 -1760 -4195 -1635
rect -4415 -2080 -4195 -1955
rect -4505 -2275 -4415 -2240
rect -5325 -2315 -5185 -2305
rect -5325 -2335 -5315 -2315
rect -5195 -2335 -5185 -2315
rect -3830 -2315 -3695 -2305
rect -3830 -2320 -3820 -2315
rect -5325 -2345 -5185 -2335
rect -4770 -2355 -3820 -2320
rect -4770 -2400 -4740 -2355
rect -3830 -2360 -3820 -2355
rect -3705 -2360 -3695 -2315
rect -3830 -2370 -3695 -2360
rect -4860 -2435 -4735 -2400
rect -10150 -2565 -9930 -2435
rect -5080 -2730 -4860 -2600
rect -4735 -2730 -4515 -2600
rect -10150 -2895 -9930 -2765
rect -3615 -2830 -3575 -1035
rect -2005 -1280 -1785 -1155
rect -2005 -1600 -1785 -1475
rect -1765 -1545 -1745 -880
rect -1690 -1245 -1670 -860
rect 245 -1020 1000 -1010
rect 245 -1040 255 -1020
rect 525 -1040 660 -1020
rect 930 -1040 1000 -1020
rect 245 -1050 1000 -1040
rect 245 -1085 535 -1075
rect 245 -1105 255 -1085
rect 525 -1105 535 -1085
rect 245 -1115 535 -1105
rect 650 -1085 940 -1075
rect 650 -1105 660 -1085
rect 930 -1105 940 -1085
rect 650 -1135 940 -1105
rect 650 -1155 660 -1135
rect 930 -1155 940 -1135
rect 650 -1195 940 -1155
rect -25 -1230 940 -1195
rect -1725 -1255 -1575 -1245
rect -1725 -1495 -1715 -1255
rect -1585 -1495 -1575 -1255
rect -1725 -1505 -1575 -1495
rect -1765 -1555 -1575 -1545
rect -1765 -1575 -1715 -1555
rect -2005 -1920 -1785 -1795
rect -1725 -1795 -1715 -1575
rect -1585 -1795 -1575 -1555
rect -1725 -1805 -1575 -1795
rect -2005 -2240 -1785 -2115
rect -25 -2830 10 -1230
rect 775 -2565 995 -2435
rect -5080 -2850 -4860 -2835
rect -5080 -2895 -5070 -2850
rect -4875 -2895 -4860 -2850
rect -4735 -2870 10 -2830
rect -4735 -2895 -4515 -2870
rect 775 -2895 995 -2765
<< viali >>
rect -8245 0 -8225 70
rect -8115 0 -8095 70
rect -7970 0 -7950 70
rect -7920 0 -7900 70
rect -7970 -205 -7950 -135
rect -7920 -205 -7900 -135
rect -7560 0 -7540 70
rect -4515 -15 -4495 55
rect -4465 -15 -4445 55
rect -7560 -205 -7540 -135
rect -4790 -220 -4770 -150
rect -4660 -220 -4640 -150
rect -4515 -220 -4495 -150
rect -4465 -220 -4445 -150
rect -7570 -425 -7510 -405
rect -4895 -420 -4835 -400
rect -7550 -565 -7530 -505
rect -7465 -1620 -7335 -1380
rect -4705 -1495 -4575 -1255
rect -4705 -1900 -4575 -1660
rect -4455 -525 -4395 -505
rect -1715 -525 -1655 -505
rect -3820 -2360 -3705 -2315
rect 255 -1105 525 -1085
rect 660 -1155 930 -1135
rect -1715 -1495 -1585 -1255
rect -1715 -1795 -1585 -1555
rect -5070 -2895 -4875 -2850
rect -5070 -2915 -4875 -2895
<< metal1 >>
rect -8255 70 -8215 145
rect -8255 0 -8245 70
rect -8225 0 -8215 70
rect -8255 -10 -8215 0
rect -8125 70 -8085 145
rect -7795 80 -7560 85
rect -8125 0 -8115 70
rect -8095 0 -8085 70
rect -8125 -10 -8085 0
rect -7980 70 -7455 80
rect -7980 0 -7970 70
rect -7950 0 -7920 70
rect -7900 0 -7560 70
rect -7540 0 -7455 70
rect -4800 55 -4385 65
rect -7980 -10 -7455 0
rect -7980 -25 -7935 -10
rect -10150 -110 -7935 -25
rect -7355 -75 -7315 15
rect -4945 -15 -4515 55
rect -4495 -15 -4465 55
rect -4445 -15 -4385 55
rect -4945 -25 -4385 -15
rect -4275 -75 -4235 -50
rect -7570 -110 -7315 -75
rect -4800 -95 -4235 -75
rect -4800 -100 -4435 -95
rect -7570 -125 -7530 -110
rect -10150 -135 -7530 -125
rect -10150 -205 -7970 -135
rect -7950 -205 -7920 -135
rect -7900 -205 -7560 -135
rect -7540 -205 -7530 -135
rect -10150 -215 -7530 -205
rect -4800 -140 -4755 -100
rect -4475 -140 -4435 -100
rect -4800 -150 -4760 -140
rect -4800 -220 -4790 -150
rect -4770 -220 -4760 -150
rect -4800 -230 -4760 -220
rect -4670 -150 -4630 -140
rect -4670 -220 -4660 -150
rect -4640 -220 -4630 -150
rect -4670 -390 -4630 -220
rect -4525 -150 -4435 -140
rect -4525 -220 -4515 -150
rect -4495 -220 -4465 -150
rect -4445 -220 -4435 -150
rect -4525 -230 -4435 -220
rect -4410 -350 -4405 -210
rect -1795 -350 -1665 -210
rect -7580 -405 -7385 -395
rect -7580 -470 -7570 -405
rect -7395 -470 -7385 -405
rect -4905 -400 -4630 -390
rect -4905 -420 -4895 -400
rect -4835 -420 -4630 -400
rect -4905 -430 -4630 -420
rect -4465 -400 -4385 -390
rect -7580 -480 -7385 -470
rect -4595 -455 -4515 -445
rect -7560 -505 -7470 -495
rect -7560 -565 -7550 -505
rect -7530 -515 -7470 -505
rect -7530 -565 -7520 -515
rect -4595 -525 -4585 -455
rect -4525 -495 -4515 -455
rect -4465 -470 -4455 -400
rect -4395 -470 -4385 -400
rect -4465 -480 -4385 -470
rect -1725 -400 -1645 -390
rect -1725 -470 -1715 -400
rect -1655 -470 -1645 -400
rect -1725 -480 -1645 -470
rect -4525 -505 -4385 -495
rect -4525 -525 -4455 -505
rect -4395 -525 -4385 -505
rect -4595 -535 -4385 -525
rect -1725 -505 -1645 -495
rect -1725 -525 -1715 -505
rect -1655 -525 -1645 -505
rect -1725 -535 -1645 -525
rect -7560 -575 -7520 -565
rect -4870 -720 -4400 -580
rect -1790 -720 -1660 -580
rect -7470 -1035 -7455 -895
rect 285 -945 375 -940
rect 245 -1005 335 -945
rect -7465 -1115 -7425 -1035
rect 245 -1085 535 -1005
rect 245 -1105 255 -1085
rect 525 -1105 535 -1085
rect 245 -1115 535 -1105
rect -7545 -1125 -7405 -1115
rect -7545 -1205 -7535 -1125
rect -7595 -1245 -7535 -1205
rect -7415 -1245 -7405 -1125
rect 650 -1135 940 -1075
rect 650 -1155 660 -1135
rect 930 -1155 940 -1135
rect 650 -1165 940 -1155
rect -7595 -1255 -7405 -1245
rect -4715 -1255 -4565 -1245
rect -7595 -2345 -7565 -1255
rect -7475 -1380 -7325 -1370
rect -7475 -1620 -7465 -1380
rect -7335 -1620 -7325 -1380
rect -4715 -1495 -4705 -1255
rect -4575 -1495 -4565 -1255
rect -4715 -1505 -4565 -1495
rect -1725 -1255 -1575 -1245
rect -1725 -1495 -1715 -1255
rect -1585 -1495 -1575 -1255
rect -1725 -1505 -1575 -1495
rect -7475 -1630 -7325 -1620
rect -1725 -1555 -1575 -1545
rect -4715 -1660 -4565 -1650
rect -4715 -1900 -4705 -1660
rect -4575 -1900 -4565 -1660
rect -1725 -1795 -1715 -1555
rect -1585 -1795 -1575 -1555
rect -1725 -1805 -1575 -1795
rect -4715 -1910 -4565 -1900
rect -5330 -2345 -5180 -2300
rect -7595 -2375 -5180 -2345
rect -3830 -2315 -3695 -2305
rect -3830 -2360 -3820 -2315
rect -3705 -2360 -3695 -2315
rect -3830 -2370 -3695 -2360
rect -5270 -2835 -5180 -2375
rect -5270 -2850 -4860 -2835
rect -5270 -2870 -5070 -2850
rect -5080 -2915 -5070 -2870
rect -4875 -2915 -4860 -2850
rect -5080 -2930 -4860 -2915
<< via1 >>
rect -7570 -425 -7510 -405
rect -7510 -425 -7395 -405
rect -7570 -470 -7395 -425
rect -4585 -525 -4525 -455
rect -4455 -470 -4395 -400
rect -1715 -470 -1655 -400
rect -7535 -1245 -7415 -1125
rect -7465 -1620 -7335 -1380
rect -4705 -1495 -4575 -1255
rect -1715 -1495 -1585 -1255
rect -4705 -1900 -4575 -1660
rect -1715 -1795 -1585 -1555
rect -3820 -2360 -3705 -2315
<< metal2 >>
rect -4460 -310 -4430 145
rect -4545 -340 -4430 -310
rect -7580 -405 -7385 -395
rect -7580 -470 -7570 -405
rect -7395 -470 -7385 -405
rect -4545 -445 -4515 -340
rect -7580 -480 -7385 -470
rect -4595 -455 -4515 -445
rect -4595 -525 -4585 -455
rect -4525 -525 -4515 -455
rect -4465 -400 -4385 -390
rect -4465 -470 -4455 -400
rect -4395 -470 -4385 -400
rect -4465 -480 -4385 -470
rect -4595 -535 -4515 -525
rect -4415 -1065 -4385 -480
rect -1725 -400 -1645 -390
rect -1725 -470 -1715 -400
rect -1655 -470 -1645 -400
rect -1725 -480 -1645 -470
rect -1725 -1060 -1695 -480
rect -2385 -1065 -1695 -1060
rect -4415 -1085 -1695 -1065
rect -7545 -1125 -7405 -1115
rect -7545 -1245 -7535 -1125
rect -7415 -1245 -7405 -1125
rect -7545 -1255 -7405 -1245
rect -4715 -1255 -4565 -1245
rect -7475 -1380 -7325 -1370
rect -7475 -1620 -7465 -1380
rect -7335 -1620 -7325 -1380
rect -4715 -1495 -4705 -1255
rect -4575 -1495 -4565 -1255
rect -4715 -1505 -4565 -1495
rect -7475 -1630 -7325 -1620
rect -4715 -1660 -4565 -1650
rect -4715 -1900 -4705 -1660
rect -4575 -1900 -4565 -1660
rect -4715 -1910 -4565 -1900
rect -2160 -2305 -2125 -1085
rect -1725 -1255 -1575 -1245
rect -1725 -1495 -1715 -1255
rect -1585 -1495 -1575 -1255
rect -1725 -1505 -1575 -1495
rect -1725 -1555 -1575 -1545
rect -1725 -1795 -1715 -1555
rect -1585 -1795 -1575 -1555
rect -1725 -1805 -1575 -1795
rect -3830 -2315 -2125 -2305
rect -3830 -2360 -3820 -2315
rect -3705 -2360 -2125 -2315
rect -3830 -2370 -2125 -2360
<< via2 >>
rect -7570 -470 -7395 -405
rect -7535 -1245 -7415 -1125
rect -7465 -1620 -7335 -1380
rect -4705 -1495 -4575 -1255
rect -4705 -1900 -4575 -1660
rect -1715 -1495 -1585 -1255
rect -1715 -1795 -1585 -1555
<< metal3 >>
rect -10150 -1115 -7620 -245
rect -7580 -405 -7385 -395
rect -7580 -470 -7570 -405
rect -7395 -470 -7385 -405
rect -7580 -480 -7385 -470
rect -10150 -1125 -7405 -1115
rect -10150 -1245 -7535 -1125
rect -7415 -1245 -7405 -1125
rect -10150 -1255 -7405 -1245
rect -7285 -1255 -4565 -1245
rect -10150 -2275 -7620 -1255
rect -7475 -1380 -7325 -1370
rect -7475 -1620 -7465 -1380
rect -7335 -1620 -7325 -1380
rect -7475 -1630 -7325 -1620
rect -7285 -1495 -4705 -1255
rect -4575 -1495 -4565 -1255
rect -7285 -1505 -4565 -1495
rect -1725 -1255 995 -1245
rect -1725 -1495 -1715 -1255
rect -1585 -1495 995 -1255
rect -1725 -1505 995 -1495
rect -7285 -2275 -4755 -1505
rect -1725 -1555 -1575 -1545
rect -4715 -1660 -4565 -1650
rect -4715 -1900 -4705 -1660
rect -4575 -1900 -4565 -1660
rect -1725 -1795 -1715 -1555
rect -1585 -1795 -1575 -1555
rect -1725 -1805 -1575 -1795
rect -4715 -1910 -4565 -1900
rect -1535 -2275 995 -1505
<< via3 >>
rect -7570 -470 -7395 -405
rect -7465 -1620 -7335 -1380
rect -4705 -1900 -4575 -1660
rect -1715 -1795 -1585 -1555
<< mimcap >>
rect -10135 -270 -7635 -260
rect -10135 -510 -7785 -270
rect -7645 -510 -7635 -270
rect -10135 -2260 -7635 -510
rect -7270 -1380 -4770 -1260
rect -7270 -1620 -7260 -1380
rect -7130 -1620 -4770 -1380
rect -7270 -1660 -4770 -1620
rect -7270 -1900 -4910 -1660
rect -4780 -1900 -4770 -1660
rect -7270 -2260 -4770 -1900
rect -1520 -1555 980 -1260
rect -1520 -1795 -1510 -1555
rect -1380 -1795 980 -1555
rect -1520 -2260 980 -1795
<< mimcapcontact >>
rect -7785 -510 -7645 -270
rect -7260 -1620 -7130 -1380
rect -4910 -1900 -4780 -1660
rect -1510 -1795 -1380 -1555
<< metal4 >>
rect -7795 -270 -7635 -260
rect -7795 -510 -7785 -270
rect -7645 -395 -7635 -270
rect -7645 -405 -7385 -395
rect -7645 -470 -7570 -405
rect -7395 -470 -7385 -405
rect -7645 -480 -7385 -470
rect -7645 -510 -7635 -480
rect -7795 -520 -7635 -510
rect -7475 -1380 -7120 -1370
rect -7475 -1620 -7465 -1380
rect -7335 -1620 -7260 -1380
rect -7130 -1620 -7120 -1380
rect -7475 -1630 -7120 -1620
rect -1725 -1555 -1370 -1545
rect -4920 -1660 -4565 -1650
rect -4920 -1900 -4910 -1660
rect -4780 -1900 -4705 -1660
rect -4575 -1900 -4565 -1660
rect -1725 -1795 -1715 -1555
rect -1585 -1795 -1510 -1555
rect -1380 -1795 -1370 -1555
rect -1725 -1805 -1370 -1795
rect -4920 -1910 -4565 -1900
use amux  amux_0
timestamp 1620340807
transform 1 0 -8210 0 1 -240
box -70 5 345 380
use sbc2  sbc2_2
timestamp 1620340936
transform 1 0 -7410 0 1 -515
box -80 -540 2585 645
use amux  amux_1
timestamp 1620340807
transform 1 0 -4755 0 1 -255
box -70 5 345 380
use sbc2  sbc2_1
timestamp 1620340936
transform 1 0 -4330 0 1 -515
box -80 -540 2585 645
use sbc2  sbc2_0
timestamp 1620340936
transform 1 0 -1590 0 1 -515
box -80 -540 2585 645
<< labels >>
rlabel metal1 -8105 145 -8105 145 1 VL
rlabel metal1 -8235 145 -8235 145 1 VH
rlabel locali -7830 145 -7830 145 1 source
rlabel poly -7585 145 -7585 145 1 samp
rlabel poly -4540 145 -4540 145 1 intc
rlabel metal2 -4445 145 -4445 145 1 OCC1
rlabel locali -1755 145 -1755 145 1 OCC2
rlabel locali 1000 -1030 1000 -1030 3 Vtrip
rlabel metal1 -10150 -170 -10150 -170 7 VN
rlabel metal1 -10150 -70 -10150 -70 7 VP
<< end >>
