magic
tech sky130A
timestamp 1620340936
<< nwell >>
rect -80 140 2570 630
<< nmos >>
rect -10 -210 50 -60
rect 100 -210 160 -60
rect 210 -210 270 -60
rect 320 -210 380 -60
rect 430 -210 490 -60
rect 540 -210 600 -60
rect 650 -210 710 -60
rect 760 -210 820 -60
rect 970 -210 1030 -60
rect 1080 -210 1140 -60
rect 1190 -210 1250 -60
rect 1300 -210 1360 -60
rect 1410 -210 1470 -60
rect 1520 -210 1580 -60
rect 1730 -210 1790 -60
rect 1840 -210 1900 -60
rect 2030 -210 2090 -60
rect 2140 -210 2200 -60
rect 2330 -210 2390 -60
rect 2440 -210 2500 -60
rect -10 -525 50 -375
rect 100 -525 160 -375
rect 210 -525 270 -375
rect 320 -525 380 -375
rect 430 -525 490 -375
rect 540 -525 600 -375
rect 650 -525 710 -375
rect 760 -525 820 -375
rect 870 -525 930 -375
rect 980 -525 1040 -375
rect 1090 -525 1150 -375
rect 1200 -525 1260 -375
rect 1310 -525 1370 -375
rect 1420 -525 1480 -375
rect 1530 -525 1590 -375
rect 1640 -525 1700 -375
rect 1835 -385 2435 -370
<< pmos >>
rect -10 460 50 610
rect 100 460 160 610
rect 210 460 270 610
rect 320 460 380 610
rect 430 460 490 610
rect 540 460 600 610
rect 650 460 710 610
rect 760 460 820 610
rect 870 460 930 610
rect 980 460 1040 610
rect 1090 460 1150 610
rect 1200 460 1260 610
rect 1310 460 1370 610
rect 1420 460 1480 610
rect 1530 460 1590 610
rect 1640 460 1700 610
rect 1870 510 2470 525
rect 1870 445 2470 460
rect -10 160 50 310
rect 100 160 160 310
rect 210 160 270 310
rect 320 160 380 310
rect 430 160 490 310
rect 540 160 600 310
rect 650 160 710 310
rect 760 160 820 310
rect 970 160 1030 310
rect 1080 160 1140 310
rect 1190 160 1250 310
rect 1300 160 1360 310
rect 1410 160 1470 310
rect 1520 160 1580 310
rect 1730 160 1790 310
rect 1840 160 1900 310
rect 2030 160 2090 310
rect 2140 160 2200 310
rect 2330 160 2390 310
rect 2440 160 2500 310
<< ndiff >>
rect -60 -75 -10 -60
rect -60 -195 -45 -75
rect -25 -195 -10 -75
rect -60 -210 -10 -195
rect 50 -75 100 -60
rect 50 -195 65 -75
rect 85 -195 100 -75
rect 50 -210 100 -195
rect 160 -75 210 -60
rect 160 -195 175 -75
rect 195 -195 210 -75
rect 160 -210 210 -195
rect 270 -75 320 -60
rect 270 -195 285 -75
rect 305 -195 320 -75
rect 270 -210 320 -195
rect 380 -75 430 -60
rect 380 -195 395 -75
rect 415 -195 430 -75
rect 380 -210 430 -195
rect 490 -75 540 -60
rect 490 -195 505 -75
rect 525 -195 540 -75
rect 490 -210 540 -195
rect 600 -75 650 -60
rect 600 -195 615 -75
rect 635 -195 650 -75
rect 600 -210 650 -195
rect 710 -75 760 -60
rect 710 -195 725 -75
rect 745 -195 760 -75
rect 710 -210 760 -195
rect 820 -75 870 -60
rect 920 -75 970 -60
rect 820 -195 835 -75
rect 855 -195 870 -75
rect 920 -195 935 -75
rect 955 -195 970 -75
rect 820 -210 870 -195
rect 920 -210 970 -195
rect 1030 -75 1080 -60
rect 1030 -195 1045 -75
rect 1065 -195 1080 -75
rect 1030 -210 1080 -195
rect 1140 -75 1190 -60
rect 1140 -195 1155 -75
rect 1175 -195 1190 -75
rect 1140 -210 1190 -195
rect 1250 -75 1300 -60
rect 1250 -195 1265 -75
rect 1285 -195 1300 -75
rect 1250 -210 1300 -195
rect 1360 -75 1410 -60
rect 1360 -195 1375 -75
rect 1395 -195 1410 -75
rect 1360 -210 1410 -195
rect 1470 -75 1520 -60
rect 1470 -195 1485 -75
rect 1505 -195 1520 -75
rect 1470 -210 1520 -195
rect 1580 -75 1630 -60
rect 1580 -195 1595 -75
rect 1615 -195 1630 -75
rect 1580 -210 1630 -195
rect 1680 -75 1730 -60
rect 1680 -195 1695 -75
rect 1715 -195 1730 -75
rect 1680 -210 1730 -195
rect 1790 -75 1840 -60
rect 1790 -195 1805 -75
rect 1825 -195 1840 -75
rect 1790 -210 1840 -195
rect 1900 -75 1950 -60
rect 1900 -195 1915 -75
rect 1935 -195 1950 -75
rect 1900 -210 1950 -195
rect 1980 -75 2030 -60
rect 1980 -195 1995 -75
rect 2015 -195 2030 -75
rect 1980 -210 2030 -195
rect 2090 -75 2140 -60
rect 2090 -195 2105 -75
rect 2125 -195 2140 -75
rect 2090 -210 2140 -195
rect 2200 -75 2250 -60
rect 2200 -195 2215 -75
rect 2235 -195 2250 -75
rect 2200 -210 2250 -195
rect 2280 -75 2330 -60
rect 2280 -195 2295 -75
rect 2315 -195 2330 -75
rect 2280 -210 2330 -195
rect 2390 -75 2440 -60
rect 2390 -195 2405 -75
rect 2425 -195 2440 -75
rect 2390 -210 2440 -195
rect 2500 -75 2550 -60
rect 2500 -195 2515 -75
rect 2535 -195 2550 -75
rect 2500 -210 2550 -195
rect 1835 -335 2435 -320
rect 1835 -355 1850 -335
rect 2420 -355 2435 -335
rect 1835 -370 2435 -355
rect -60 -390 -10 -375
rect -60 -510 -45 -390
rect -25 -510 -10 -390
rect -60 -525 -10 -510
rect 50 -390 100 -375
rect 50 -510 65 -390
rect 85 -510 100 -390
rect 50 -525 100 -510
rect 160 -390 210 -375
rect 160 -510 175 -390
rect 195 -510 210 -390
rect 160 -525 210 -510
rect 270 -390 320 -375
rect 270 -510 285 -390
rect 305 -510 320 -390
rect 270 -525 320 -510
rect 380 -390 430 -375
rect 380 -510 395 -390
rect 415 -510 430 -390
rect 380 -525 430 -510
rect 490 -390 540 -375
rect 490 -510 505 -390
rect 525 -510 540 -390
rect 490 -525 540 -510
rect 600 -390 650 -375
rect 600 -510 615 -390
rect 635 -510 650 -390
rect 600 -525 650 -510
rect 710 -390 760 -375
rect 710 -510 725 -390
rect 745 -510 760 -390
rect 710 -525 760 -510
rect 820 -390 870 -375
rect 820 -510 835 -390
rect 855 -510 870 -390
rect 820 -525 870 -510
rect 930 -390 980 -375
rect 930 -510 945 -390
rect 965 -510 980 -390
rect 930 -525 980 -510
rect 1040 -390 1090 -375
rect 1040 -510 1055 -390
rect 1075 -510 1090 -390
rect 1040 -525 1090 -510
rect 1150 -390 1200 -375
rect 1150 -510 1165 -390
rect 1185 -510 1200 -390
rect 1150 -525 1200 -510
rect 1260 -390 1310 -375
rect 1260 -510 1275 -390
rect 1295 -510 1310 -390
rect 1260 -525 1310 -510
rect 1370 -390 1420 -375
rect 1370 -510 1385 -390
rect 1405 -510 1420 -390
rect 1370 -525 1420 -510
rect 1480 -390 1530 -375
rect 1480 -510 1495 -390
rect 1515 -510 1530 -390
rect 1480 -525 1530 -510
rect 1590 -390 1640 -375
rect 1590 -510 1605 -390
rect 1625 -510 1640 -390
rect 1590 -525 1640 -510
rect 1700 -390 1750 -375
rect 1700 -510 1715 -390
rect 1735 -510 1750 -390
rect 1835 -400 2435 -385
rect 1835 -420 1850 -400
rect 2420 -420 2435 -400
rect 1835 -435 2435 -420
rect 1700 -525 1750 -510
<< pdiff >>
rect -60 595 -10 610
rect -60 475 -45 595
rect -25 475 -10 595
rect -60 460 -10 475
rect 50 595 100 610
rect 50 475 65 595
rect 85 475 100 595
rect 50 460 100 475
rect 160 595 210 610
rect 160 475 175 595
rect 195 475 210 595
rect 160 460 210 475
rect 270 595 320 610
rect 270 475 285 595
rect 305 475 320 595
rect 270 460 320 475
rect 380 595 430 610
rect 380 475 395 595
rect 415 475 430 595
rect 380 460 430 475
rect 490 595 540 610
rect 490 475 505 595
rect 525 475 540 595
rect 490 460 540 475
rect 600 595 650 610
rect 600 475 615 595
rect 635 475 650 595
rect 600 460 650 475
rect 710 595 760 610
rect 710 475 725 595
rect 745 475 760 595
rect 710 460 760 475
rect 820 595 870 610
rect 820 475 835 595
rect 855 475 870 595
rect 820 460 870 475
rect 930 595 980 610
rect 930 475 945 595
rect 965 475 980 595
rect 930 460 980 475
rect 1040 595 1090 610
rect 1040 475 1055 595
rect 1075 475 1090 595
rect 1040 460 1090 475
rect 1150 595 1200 610
rect 1150 475 1165 595
rect 1185 475 1200 595
rect 1150 460 1200 475
rect 1260 595 1310 610
rect 1260 475 1275 595
rect 1295 475 1310 595
rect 1260 460 1310 475
rect 1370 595 1420 610
rect 1370 475 1385 595
rect 1405 475 1420 595
rect 1370 460 1420 475
rect 1480 595 1530 610
rect 1480 475 1495 595
rect 1515 475 1530 595
rect 1480 460 1530 475
rect 1590 595 1640 610
rect 1590 475 1605 595
rect 1625 475 1640 595
rect 1590 460 1640 475
rect 1700 595 1750 610
rect 1700 475 1715 595
rect 1735 475 1750 595
rect 1870 560 2470 575
rect 1870 540 1885 560
rect 2455 540 2470 560
rect 1870 525 2470 540
rect 1700 460 1750 475
rect 1870 495 2470 510
rect 1870 475 1885 495
rect 2455 475 2470 495
rect 1870 460 2470 475
rect 1870 430 2470 445
rect 1870 410 1885 430
rect 2455 410 2470 430
rect 1870 395 2470 410
rect -60 295 -10 310
rect -60 175 -45 295
rect -25 175 -10 295
rect -60 160 -10 175
rect 50 295 100 310
rect 50 175 65 295
rect 85 175 100 295
rect 50 160 100 175
rect 160 295 210 310
rect 160 175 175 295
rect 195 175 210 295
rect 160 160 210 175
rect 270 295 320 310
rect 270 175 285 295
rect 305 175 320 295
rect 270 160 320 175
rect 380 295 430 310
rect 380 175 395 295
rect 415 175 430 295
rect 380 160 430 175
rect 490 295 540 310
rect 490 175 505 295
rect 525 175 540 295
rect 490 160 540 175
rect 600 295 650 310
rect 600 175 615 295
rect 635 175 650 295
rect 600 160 650 175
rect 710 295 760 310
rect 710 175 725 295
rect 745 175 760 295
rect 710 160 760 175
rect 820 295 870 310
rect 920 295 970 310
rect 820 175 835 295
rect 855 175 870 295
rect 920 175 935 295
rect 955 175 970 295
rect 820 160 870 175
rect 920 160 970 175
rect 1030 295 1080 310
rect 1030 175 1045 295
rect 1065 175 1080 295
rect 1030 160 1080 175
rect 1140 295 1190 310
rect 1140 175 1155 295
rect 1175 175 1190 295
rect 1140 160 1190 175
rect 1250 295 1300 310
rect 1250 175 1265 295
rect 1285 175 1300 295
rect 1250 160 1300 175
rect 1360 295 1410 310
rect 1360 175 1375 295
rect 1395 175 1410 295
rect 1360 160 1410 175
rect 1470 295 1520 310
rect 1470 175 1485 295
rect 1505 175 1520 295
rect 1470 160 1520 175
rect 1580 295 1630 310
rect 1580 175 1595 295
rect 1615 175 1630 295
rect 1580 160 1630 175
rect 1680 295 1730 310
rect 1680 175 1695 295
rect 1715 175 1730 295
rect 1680 160 1730 175
rect 1790 295 1840 310
rect 1790 175 1805 295
rect 1825 175 1840 295
rect 1790 160 1840 175
rect 1900 295 1950 310
rect 1900 175 1915 295
rect 1935 175 1950 295
rect 1900 160 1950 175
rect 1980 295 2030 310
rect 1980 175 1995 295
rect 2015 175 2030 295
rect 1980 160 2030 175
rect 2090 295 2140 310
rect 2090 175 2105 295
rect 2125 175 2140 295
rect 2090 160 2140 175
rect 2200 295 2250 310
rect 2200 175 2215 295
rect 2235 175 2250 295
rect 2200 160 2250 175
rect 2280 295 2330 310
rect 2280 175 2295 295
rect 2315 175 2330 295
rect 2280 160 2330 175
rect 2390 295 2440 310
rect 2390 175 2405 295
rect 2425 175 2440 295
rect 2390 160 2440 175
rect 2500 295 2550 310
rect 2500 175 2515 295
rect 2535 175 2550 295
rect 2500 160 2550 175
<< ndiffc >>
rect -45 -195 -25 -75
rect 65 -195 85 -75
rect 175 -195 195 -75
rect 285 -195 305 -75
rect 395 -195 415 -75
rect 505 -195 525 -75
rect 615 -195 635 -75
rect 725 -195 745 -75
rect 835 -195 855 -75
rect 935 -195 955 -75
rect 1045 -195 1065 -75
rect 1155 -195 1175 -75
rect 1265 -195 1285 -75
rect 1375 -195 1395 -75
rect 1485 -195 1505 -75
rect 1595 -195 1615 -75
rect 1695 -195 1715 -75
rect 1805 -195 1825 -75
rect 1915 -195 1935 -75
rect 1995 -195 2015 -75
rect 2105 -195 2125 -75
rect 2215 -195 2235 -75
rect 2295 -195 2315 -75
rect 2405 -195 2425 -75
rect 2515 -195 2535 -75
rect 1850 -355 2420 -335
rect -45 -510 -25 -390
rect 65 -510 85 -390
rect 175 -510 195 -390
rect 285 -510 305 -390
rect 395 -510 415 -390
rect 505 -510 525 -390
rect 615 -510 635 -390
rect 725 -510 745 -390
rect 835 -510 855 -390
rect 945 -510 965 -390
rect 1055 -510 1075 -390
rect 1165 -510 1185 -390
rect 1275 -510 1295 -390
rect 1385 -510 1405 -390
rect 1495 -510 1515 -390
rect 1605 -510 1625 -390
rect 1715 -510 1735 -390
rect 1850 -420 2420 -400
<< pdiffc >>
rect -45 475 -25 595
rect 65 475 85 595
rect 175 475 195 595
rect 285 475 305 595
rect 395 475 415 595
rect 505 475 525 595
rect 615 475 635 595
rect 725 475 745 595
rect 835 475 855 595
rect 945 475 965 595
rect 1055 475 1075 595
rect 1165 475 1185 595
rect 1275 475 1295 595
rect 1385 475 1405 595
rect 1495 475 1515 595
rect 1605 475 1625 595
rect 1715 475 1735 595
rect 1885 540 2455 560
rect 1885 475 2455 495
rect 1885 410 2455 430
rect -45 175 -25 295
rect 65 175 85 295
rect 175 175 195 295
rect 285 175 305 295
rect 395 175 415 295
rect 505 175 525 295
rect 615 175 635 295
rect 725 175 745 295
rect 835 175 855 295
rect 935 175 955 295
rect 1045 175 1065 295
rect 1155 175 1175 295
rect 1265 175 1285 295
rect 1375 175 1395 295
rect 1485 175 1505 295
rect 1595 175 1615 295
rect 1695 175 1715 295
rect 1805 175 1825 295
rect 1915 175 1935 295
rect 1995 175 2015 295
rect 2105 175 2125 295
rect 2215 175 2235 295
rect 2295 175 2315 295
rect 2405 175 2425 295
rect 2515 175 2535 295
<< psubdiff >>
rect 870 -75 920 -60
rect 870 -195 885 -75
rect 905 -195 920 -75
rect 870 -210 920 -195
rect 1750 -390 1800 -375
rect 1750 -510 1765 -390
rect 1785 -510 1800 -390
rect 1750 -525 1800 -510
<< nsubdiff >>
rect 1750 595 1800 610
rect 1750 475 1765 595
rect 1785 475 1800 595
rect 1750 460 1800 475
rect 870 295 920 310
rect 870 175 885 295
rect 905 175 920 295
rect 870 160 920 175
<< psubdiffcont >>
rect 885 -195 905 -75
rect 1765 -510 1785 -390
<< nsubdiffcont >>
rect 1765 475 1785 595
rect 885 175 905 295
<< poly >>
rect -10 610 50 625
rect 100 620 710 635
rect 100 610 160 620
rect 210 610 270 620
rect 320 610 380 620
rect 430 610 490 620
rect 540 610 600 620
rect 650 610 710 620
rect 760 610 820 625
rect 870 610 930 625
rect 980 620 1590 635
rect 980 610 1040 620
rect 1090 610 1150 620
rect 1200 610 1260 620
rect 1310 610 1370 620
rect 1420 610 1480 620
rect 1530 610 1590 620
rect 1640 610 1700 625
rect 1810 510 1870 525
rect 2470 510 2495 525
rect 1810 460 1860 510
rect 2480 460 2495 510
rect -10 445 50 460
rect 100 445 160 460
rect 210 445 270 460
rect 320 445 380 460
rect 430 445 490 460
rect 540 445 600 460
rect 650 445 710 460
rect -10 435 30 445
rect -10 415 0 435
rect 20 415 30 435
rect -10 405 30 415
rect -10 355 30 365
rect -10 335 0 355
rect 20 335 30 355
rect 145 335 160 445
rect 255 335 270 445
rect 365 335 380 445
rect 475 335 490 445
rect 585 335 600 445
rect 695 405 710 445
rect 760 450 820 460
rect 870 450 930 460
rect 760 435 930 450
rect 890 415 900 435
rect 920 415 930 435
rect 890 405 930 415
rect 980 450 1040 460
rect 1090 450 1150 460
rect 980 435 1150 450
rect 1200 445 1260 460
rect 1310 445 1370 460
rect 1420 445 1480 460
rect 1530 445 1590 460
rect 1640 435 1700 460
rect 695 390 860 405
rect 695 335 710 390
rect 845 375 860 390
rect 980 375 995 435
rect 1045 415 1055 435
rect 1075 415 1085 435
rect 1045 405 1085 415
rect 1640 415 1670 435
rect 1690 415 1700 435
rect 1640 405 1700 415
rect 1810 445 1870 460
rect 2470 445 2495 460
rect 1810 405 1860 445
rect -10 325 30 335
rect -10 310 50 325
rect 100 320 710 335
rect 780 355 820 365
rect 845 360 995 375
rect 1125 360 1425 375
rect 780 335 790 355
rect 810 335 820 355
rect 780 325 1030 335
rect 1125 325 1140 360
rect 100 310 160 320
rect 210 310 270 320
rect 320 310 380 320
rect 430 310 490 320
rect 540 310 600 320
rect 650 310 710 320
rect 760 320 1030 325
rect 760 310 820 320
rect 970 310 1030 320
rect 1080 310 1140 325
rect 1190 320 1360 335
rect 1190 310 1250 320
rect 1300 310 1360 320
rect 1410 325 1425 360
rect 1640 335 1660 405
rect 1790 395 1860 405
rect 1790 375 1800 395
rect 1820 375 1860 395
rect 1790 365 1860 375
rect 2460 355 2500 365
rect 2460 335 2470 355
rect 2490 335 2500 355
rect 1410 310 1470 325
rect 1520 320 1790 335
rect 2460 325 2500 335
rect 1520 310 1580 320
rect 1730 310 1790 320
rect 1840 310 1900 325
rect 2030 310 2090 325
rect 2140 310 2200 325
rect 2330 310 2390 325
rect 2440 310 2500 325
rect -10 145 50 160
rect 100 145 160 160
rect 210 145 270 160
rect 320 145 380 160
rect 430 145 490 160
rect 540 145 600 160
rect 650 145 710 160
rect 760 145 820 160
rect 970 145 1030 160
rect 1080 145 1140 160
rect 1190 145 1250 160
rect 1300 145 1360 160
rect 1410 145 1470 160
rect 1520 150 1580 160
rect 1730 150 1790 160
rect 115 105 155 115
rect 115 85 125 105
rect 145 85 155 105
rect 115 75 155 85
rect -10 -20 30 -10
rect -10 -40 0 -20
rect 20 -40 30 -20
rect 115 -35 130 75
rect 695 30 710 145
rect 1190 100 1225 145
rect 1410 100 1445 145
rect 1520 135 1790 150
rect 1840 150 1900 160
rect 2030 150 2090 160
rect 2140 150 2200 160
rect 2330 150 2390 160
rect 1840 135 2390 150
rect 2440 145 2500 160
rect 1100 50 1225 100
rect 1320 60 1445 100
rect 1100 30 1140 50
rect 695 20 750 30
rect 695 0 720 20
rect 740 0 750 20
rect 695 -10 750 0
rect 1100 10 1110 30
rect 1130 10 1140 30
rect 780 -20 820 -10
rect -10 -45 30 -40
rect -10 -60 50 -45
rect 100 -50 710 -35
rect 780 -40 790 -20
rect 810 -35 820 -20
rect 810 -40 1030 -35
rect 780 -45 1030 -40
rect 1100 -45 1140 10
rect 1320 30 1360 60
rect 1320 10 1330 30
rect 1350 10 1360 30
rect 1320 -35 1360 10
rect 1860 -10 1900 135
rect 2330 -10 2370 135
rect 1540 -20 1580 -10
rect 1540 -35 1550 -20
rect 100 -60 160 -50
rect 210 -60 270 -50
rect 320 -60 380 -50
rect 430 -60 490 -50
rect 540 -60 600 -50
rect 650 -60 710 -50
rect 760 -50 1030 -45
rect 760 -60 820 -50
rect 970 -60 1030 -50
rect 1080 -60 1140 -45
rect 1190 -50 1360 -35
rect 1520 -40 1550 -35
rect 1570 -35 1580 -20
rect 1730 -20 1770 -10
rect 1730 -35 1740 -20
rect 1570 -40 1740 -35
rect 1760 -35 1770 -20
rect 1860 -20 2370 -10
rect 1860 -35 1870 -20
rect 1760 -40 1790 -35
rect 1190 -60 1250 -50
rect 1300 -60 1360 -50
rect 1410 -60 1470 -45
rect 1520 -50 1790 -40
rect 1520 -60 1580 -50
rect 1730 -60 1790 -50
rect 1840 -40 1870 -35
rect 1890 -40 2340 -20
rect 2360 -35 2370 -20
rect 2460 -20 2500 -10
rect 2360 -40 2390 -35
rect 1840 -50 2390 -40
rect 2460 -40 2470 -20
rect 2490 -40 2500 -20
rect 2460 -45 2500 -40
rect 1840 -60 1900 -50
rect 2030 -60 2090 -50
rect 2140 -60 2200 -50
rect 2330 -60 2390 -50
rect 2440 -60 2500 -45
rect -10 -225 50 -210
rect 100 -225 160 -210
rect 210 -225 270 -210
rect 320 -225 380 -210
rect 430 -225 490 -210
rect 540 -225 600 -210
rect 650 -225 710 -210
rect 760 -225 820 -210
rect 970 -225 1030 -210
rect 1080 -225 1140 -210
rect 1190 -225 1250 -210
rect 1300 -225 1360 -210
rect 1410 -225 1470 -210
rect 1520 -220 1580 -210
rect 1730 -220 1790 -210
rect -10 -335 30 -325
rect -10 -355 0 -335
rect 20 -355 30 -335
rect -10 -360 30 -355
rect 100 -350 115 -225
rect 1125 -250 1140 -225
rect 1410 -250 1425 -225
rect 1520 -235 1790 -220
rect 1840 -225 1900 -210
rect 2030 -225 2090 -210
rect 2140 -225 2200 -210
rect 2225 -230 2265 -220
rect 2330 -225 2390 -210
rect 2440 -225 2500 -210
rect 1125 -265 1425 -250
rect 2225 -250 2235 -230
rect 2255 -250 2265 -230
rect 2225 -260 2465 -250
rect 2250 -275 2465 -260
rect 695 -300 865 -285
rect 695 -350 710 -300
rect 850 -310 865 -300
rect 850 -325 995 -310
rect -10 -375 50 -360
rect 100 -365 710 -350
rect 780 -335 820 -325
rect 780 -355 790 -335
rect 810 -350 820 -335
rect 980 -350 995 -325
rect 1045 -335 1085 -325
rect 1045 -350 1055 -335
rect 810 -355 930 -350
rect 780 -360 930 -355
rect 100 -375 160 -365
rect 210 -375 270 -365
rect 320 -375 380 -365
rect 430 -375 490 -365
rect 540 -375 600 -365
rect 650 -375 710 -365
rect 760 -365 930 -360
rect 760 -375 820 -365
rect 870 -375 930 -365
rect 980 -355 1055 -350
rect 1075 -350 1085 -335
rect 1660 -335 1700 -325
rect 1075 -355 1590 -350
rect 980 -365 1590 -355
rect 1660 -355 1670 -335
rect 1690 -355 1700 -335
rect 1660 -360 1700 -355
rect 980 -375 1040 -365
rect 1090 -375 1150 -365
rect 1200 -375 1260 -365
rect 1310 -375 1370 -365
rect 1420 -375 1480 -365
rect 1530 -375 1590 -365
rect 1640 -375 1700 -360
rect 2445 -365 2465 -275
rect 2445 -370 2490 -365
rect 1820 -385 1835 -370
rect 2435 -375 2490 -370
rect 2435 -385 2460 -375
rect 2450 -395 2460 -385
rect 2480 -395 2490 -375
rect 2450 -405 2490 -395
rect -10 -540 50 -525
rect 100 -540 160 -525
rect 210 -540 270 -525
rect 320 -540 380 -525
rect 430 -540 490 -525
rect 540 -540 600 -525
rect 650 -540 710 -525
rect 760 -540 820 -525
rect 870 -540 930 -525
rect 980 -540 1040 -525
rect 1090 -540 1150 -525
rect 1200 -540 1260 -525
rect 1310 -540 1370 -525
rect 1420 -540 1480 -525
rect 1530 -540 1590 -525
rect 1640 -540 1700 -525
<< polycont >>
rect 0 415 20 435
rect 0 335 20 355
rect 900 415 920 435
rect 1055 415 1075 435
rect 1670 415 1690 435
rect 790 335 810 355
rect 1800 375 1820 395
rect 2470 335 2490 355
rect 125 85 145 105
rect 0 -40 20 -20
rect 720 0 740 20
rect 1110 10 1130 30
rect 790 -40 810 -20
rect 1330 10 1350 30
rect 1550 -40 1570 -20
rect 1740 -40 1760 -20
rect 1870 -40 1890 -20
rect 2340 -40 2360 -20
rect 2470 -40 2490 -20
rect 0 -355 20 -335
rect 2235 -250 2255 -230
rect 790 -355 810 -335
rect 1055 -355 1075 -335
rect 1670 -355 1690 -335
rect 2460 -395 2480 -375
<< locali >>
rect 185 625 625 645
rect 185 605 205 625
rect -60 595 -15 605
rect -60 475 -45 595
rect -25 475 -15 595
rect -60 465 -15 475
rect 55 595 95 605
rect 55 475 65 595
rect 85 475 95 595
rect 55 465 95 475
rect 165 595 205 605
rect 165 475 175 595
rect 195 475 205 595
rect 165 465 205 475
rect 275 595 315 605
rect 275 475 285 595
rect 305 475 315 595
rect 275 465 315 475
rect 385 595 425 625
rect 605 605 625 625
rect 1155 625 1615 645
rect 1155 605 1175 625
rect 1595 605 1615 625
rect 385 475 395 595
rect 415 475 425 595
rect 385 465 425 475
rect 495 595 535 605
rect 495 475 505 595
rect 525 475 535 595
rect 495 465 535 475
rect 605 595 645 605
rect 605 475 615 595
rect 635 475 645 595
rect 605 465 645 475
rect 715 595 755 605
rect 715 475 725 595
rect 745 475 755 595
rect 715 465 755 475
rect 825 595 865 605
rect 825 475 835 595
rect 855 475 865 595
rect 825 465 865 475
rect 935 595 975 605
rect 935 475 945 595
rect 965 475 975 595
rect 935 465 975 475
rect -35 445 -15 465
rect -35 435 30 445
rect -35 425 0 435
rect -10 415 0 425
rect 20 415 30 435
rect -10 405 30 415
rect -10 355 30 365
rect -10 345 0 355
rect -35 335 0 345
rect 20 335 30 355
rect -35 325 30 335
rect 185 345 205 465
rect 845 445 865 465
rect 845 435 930 445
rect 845 425 900 435
rect 890 415 900 425
rect 920 415 930 435
rect 890 405 930 415
rect 955 365 975 465
rect 1045 595 1085 605
rect 1045 475 1055 595
rect 1075 475 1085 595
rect 1045 435 1085 475
rect 1045 415 1055 435
rect 1075 415 1085 435
rect 1045 405 1085 415
rect 1155 595 1195 605
rect 1155 475 1165 595
rect 1185 475 1195 595
rect 1155 465 1195 475
rect 1265 595 1305 605
rect 1265 475 1275 595
rect 1295 475 1305 595
rect 1265 465 1305 475
rect 1375 595 1415 605
rect 1375 475 1385 595
rect 1405 475 1415 595
rect 1375 465 1415 475
rect 1485 595 1525 605
rect 1485 475 1495 595
rect 1515 475 1525 595
rect 1485 465 1525 475
rect 1595 595 1635 605
rect 1595 475 1605 595
rect 1625 475 1635 595
rect 1595 465 1635 475
rect 1155 405 1175 465
rect 1395 445 1415 465
rect 1395 435 1560 445
rect 1395 425 1490 435
rect 1480 415 1490 425
rect 1550 415 1560 435
rect 1480 405 1560 415
rect 1120 385 1450 405
rect 1120 365 1140 385
rect 780 355 820 365
rect 185 325 625 345
rect 780 335 790 355
rect 810 345 820 355
rect 955 345 1140 365
rect 1345 355 1385 365
rect 1345 345 1355 355
rect 810 335 845 345
rect 780 325 845 335
rect -35 305 -15 325
rect 185 305 205 325
rect 605 305 625 325
rect 825 305 845 325
rect 1165 335 1355 345
rect 1375 335 1385 355
rect 1165 325 1385 335
rect 1165 305 1185 325
rect 1365 305 1385 325
rect -60 295 -15 305
rect -60 175 -45 295
rect -25 175 -15 295
rect -60 165 -15 175
rect 55 295 95 305
rect 55 175 65 295
rect 85 175 95 295
rect 55 165 95 175
rect 165 295 205 305
rect 165 175 175 295
rect 195 175 205 295
rect 165 165 205 175
rect 275 295 315 305
rect 275 175 285 295
rect 305 175 315 295
rect 275 165 315 175
rect 385 295 425 305
rect 385 175 395 295
rect 415 175 425 295
rect 385 165 425 175
rect 495 295 535 305
rect 495 175 505 295
rect 525 175 535 295
rect 495 165 535 175
rect 605 295 645 305
rect 605 175 615 295
rect 635 175 645 295
rect 605 165 645 175
rect 715 295 755 305
rect 715 175 725 295
rect 745 175 755 295
rect 715 165 755 175
rect 825 295 965 305
rect 825 175 835 295
rect 855 175 885 295
rect 905 175 935 295
rect 955 175 965 295
rect 825 165 965 175
rect 1035 295 1075 305
rect 1035 175 1045 295
rect 1065 175 1075 295
rect 1035 165 1075 175
rect 1145 295 1185 305
rect 1145 175 1155 295
rect 1175 175 1185 295
rect 1145 165 1185 175
rect 1255 295 1295 305
rect 1255 175 1265 295
rect 1285 175 1295 295
rect 1255 165 1295 175
rect 1365 295 1405 305
rect 1365 175 1375 295
rect 1395 175 1405 295
rect 1365 165 1405 175
rect 75 150 95 165
rect 75 140 155 150
rect 75 120 85 140
rect 145 120 155 140
rect 75 110 155 120
rect 115 105 155 110
rect 115 85 125 105
rect 145 85 155 105
rect 115 75 155 85
rect 405 90 425 165
rect 715 150 735 165
rect 1035 150 1055 165
rect 655 140 735 150
rect 655 120 665 140
rect 725 120 735 140
rect 655 110 735 120
rect 975 140 1055 150
rect 1255 140 1275 165
rect 975 120 985 140
rect 1045 120 1055 140
rect 975 110 1055 120
rect 1075 120 1275 140
rect 1075 90 1095 120
rect 405 70 1095 90
rect 1120 65 1200 75
rect 1120 45 1130 65
rect 1190 45 1200 65
rect 1120 40 1200 45
rect 1430 40 1450 385
rect 1475 295 1515 305
rect 1475 175 1485 295
rect 1505 175 1515 295
rect 1475 140 1515 175
rect 1475 120 1485 140
rect 1505 120 1515 140
rect 1475 110 1515 120
rect 1540 90 1560 405
rect 1615 345 1635 465
rect 1705 595 1795 605
rect 1705 475 1715 595
rect 1735 475 1765 595
rect 1785 475 1795 595
rect 1875 560 2465 570
rect 1875 540 1885 560
rect 2455 540 2465 560
rect 1875 530 2465 540
rect 1705 465 1795 475
rect 1875 495 2585 505
rect 1875 475 1885 495
rect 2455 475 2585 495
rect 1875 465 2585 475
rect 1705 445 1725 465
rect 1660 435 1725 445
rect 1660 415 1670 435
rect 1690 425 1725 435
rect 1875 430 2465 440
rect 1690 415 1700 425
rect 1660 405 1700 415
rect 1875 410 1885 430
rect 2455 410 2465 430
rect 1750 395 1830 405
rect 1875 400 2465 410
rect 1750 375 1760 395
rect 1820 375 1830 395
rect 1750 365 1830 375
rect 2460 355 2500 365
rect 1615 325 2415 345
rect 2460 335 2470 355
rect 2490 345 2500 355
rect 2490 335 2525 345
rect 2460 325 2525 335
rect 1795 305 1815 325
rect 2395 305 2415 325
rect 2505 305 2525 325
rect 1585 295 1625 305
rect 1585 175 1595 295
rect 1615 175 1625 295
rect 1585 165 1625 175
rect 1685 295 1725 305
rect 1685 175 1695 295
rect 1715 175 1725 295
rect 1685 165 1725 175
rect 1795 295 1835 305
rect 1795 175 1805 295
rect 1825 175 1835 295
rect 1795 165 1835 175
rect 1905 295 1945 305
rect 1905 175 1915 295
rect 1935 175 1945 295
rect 1905 165 1945 175
rect 1985 295 2025 305
rect 1985 175 1995 295
rect 2015 175 2025 295
rect 1985 165 2025 175
rect 2095 295 2135 305
rect 2095 175 2105 295
rect 2125 175 2135 295
rect 2095 165 2135 175
rect 2205 295 2245 305
rect 2205 175 2215 295
rect 2235 175 2245 295
rect 2205 165 2245 175
rect 2285 295 2325 305
rect 2285 175 2295 295
rect 2315 175 2325 295
rect 2285 165 2325 175
rect 2395 295 2435 305
rect 2395 175 2405 295
rect 2425 175 2435 295
rect 2395 165 2435 175
rect 2505 295 2545 305
rect 2505 175 2515 295
rect 2535 175 2545 295
rect 2505 165 2545 175
rect 1100 35 1200 40
rect 1100 30 1140 35
rect 710 20 750 30
rect 710 0 720 20
rect 740 0 750 20
rect 1100 10 1110 30
rect 1130 10 1140 30
rect 1100 0 1140 10
rect 1280 30 1360 40
rect 1280 10 1290 30
rect 1350 10 1360 30
rect 1280 0 1360 10
rect 1410 30 1450 40
rect 1410 10 1420 30
rect 1440 10 1450 30
rect 1410 0 1450 10
rect 1475 70 1560 90
rect 710 -10 750 0
rect -10 -20 30 -10
rect -10 -30 0 -20
rect -35 -40 0 -30
rect 20 -40 30 -20
rect 710 -25 735 -10
rect -35 -50 30 -40
rect 75 -45 735 -25
rect -35 -65 -15 -50
rect 75 -65 95 -45
rect 715 -65 735 -45
rect 780 -20 820 -10
rect 1475 -20 1495 70
rect 1515 40 1665 50
rect 1515 20 1525 40
rect 1585 20 1665 40
rect 1515 10 1665 20
rect 780 -40 790 -20
rect 810 -30 820 -20
rect 810 -40 845 -30
rect 780 -50 845 -40
rect 825 -65 845 -50
rect 1055 -40 1495 -20
rect 1055 -65 1075 -40
rect 1475 -65 1495 -40
rect 1540 -20 1580 -10
rect 1540 -40 1550 -20
rect 1570 -30 1580 -20
rect 1570 -40 1605 -30
rect 1540 -50 1605 -40
rect 1585 -65 1605 -50
rect -60 -75 -15 -65
rect -60 -195 -45 -75
rect -25 -195 -15 -75
rect -60 -205 -15 -195
rect 55 -75 95 -65
rect 55 -195 65 -75
rect 85 -195 95 -75
rect 55 -205 95 -195
rect 165 -75 205 -65
rect 165 -195 175 -75
rect 195 -195 205 -75
rect 165 -205 205 -195
rect 275 -75 315 -65
rect 275 -195 285 -75
rect 305 -195 315 -75
rect 275 -205 315 -195
rect 385 -75 425 -65
rect 385 -195 395 -75
rect 415 -195 425 -75
rect 385 -205 425 -195
rect 495 -75 535 -65
rect 495 -195 505 -75
rect 525 -195 535 -75
rect 495 -205 535 -195
rect 605 -75 645 -65
rect 605 -195 615 -75
rect 635 -195 645 -75
rect 605 -205 645 -195
rect 715 -75 755 -65
rect 715 -195 725 -75
rect 745 -195 755 -75
rect 715 -205 755 -195
rect 825 -75 970 -65
rect 825 -195 835 -75
rect 855 -195 885 -75
rect 905 -195 935 -75
rect 955 -195 970 -75
rect 825 -205 970 -195
rect 1035 -75 1075 -65
rect 1035 -195 1045 -75
rect 1065 -195 1075 -75
rect 1035 -205 1075 -195
rect 1145 -75 1185 -65
rect 1145 -195 1155 -75
rect 1175 -195 1185 -75
rect 1145 -205 1185 -195
rect 1255 -75 1295 -65
rect 1255 -195 1265 -75
rect 1285 -195 1295 -75
rect 1255 -205 1295 -195
rect 1365 -75 1405 -65
rect 1365 -195 1375 -75
rect 1395 -195 1405 -75
rect 1365 -205 1405 -195
rect 1475 -75 1515 -65
rect 1475 -195 1485 -75
rect 1505 -195 1515 -75
rect 1475 -205 1515 -195
rect 1585 -75 1625 -65
rect 1585 -195 1595 -75
rect 1615 -195 1625 -75
rect 1585 -205 1625 -195
rect -35 -325 -15 -205
rect 185 -225 205 -205
rect 185 -235 265 -225
rect 185 -255 195 -235
rect 255 -255 265 -235
rect 185 -265 265 -255
rect -35 -335 30 -325
rect -35 -355 0 -335
rect 20 -355 30 -335
rect -35 -365 30 -355
rect 185 -340 205 -265
rect 405 -285 425 -205
rect 605 -225 625 -205
rect 1165 -225 1185 -205
rect 1365 -225 1385 -205
rect 545 -235 625 -225
rect 545 -255 555 -235
rect 615 -255 625 -235
rect 545 -265 625 -255
rect 645 -245 1385 -225
rect 645 -285 665 -245
rect 1645 -285 1665 10
rect 1905 -10 1925 165
rect 1730 -20 1770 -10
rect 1730 -30 1740 -20
rect 1705 -40 1740 -30
rect 1760 -40 1770 -20
rect 1705 -50 1770 -40
rect 1860 -20 1925 -10
rect 1860 -40 1870 -20
rect 1890 -40 1925 -20
rect 1860 -50 1925 -40
rect 1705 -65 1725 -50
rect 1905 -65 1925 -50
rect 2005 145 2025 165
rect 2205 145 2225 165
rect 2005 125 2225 145
rect 2005 -65 2025 125
rect 2205 -65 2225 125
rect 2305 -10 2325 165
rect 2305 -20 2370 -10
rect 2305 -40 2340 -20
rect 2360 -40 2370 -20
rect 2305 -50 2370 -40
rect 2460 -20 2500 -10
rect 2460 -40 2470 -20
rect 2490 -25 2500 -20
rect 2490 -40 2525 -25
rect 2460 -50 2525 -40
rect 2305 -65 2325 -50
rect 2505 -65 2525 -50
rect 1685 -75 1725 -65
rect 1685 -195 1695 -75
rect 1715 -195 1725 -75
rect 1685 -205 1725 -195
rect 1795 -75 1835 -65
rect 1795 -195 1805 -75
rect 1825 -195 1835 -75
rect 1795 -205 1835 -195
rect 1905 -75 1945 -65
rect 1905 -195 1915 -75
rect 1935 -195 1945 -75
rect 1905 -205 1945 -195
rect 1985 -75 2025 -65
rect 1985 -195 1995 -75
rect 2015 -195 2025 -75
rect 1985 -205 2025 -195
rect 2095 -75 2135 -65
rect 2095 -195 2105 -75
rect 2125 -195 2135 -75
rect 2095 -205 2135 -195
rect 2205 -75 2245 -65
rect 2205 -195 2215 -75
rect 2235 -195 2245 -75
rect 2205 -205 2245 -195
rect 2285 -75 2325 -65
rect 2285 -195 2295 -75
rect 2315 -195 2325 -75
rect 2285 -205 2325 -195
rect 2395 -75 2435 -65
rect 2395 -195 2405 -75
rect 2425 -195 2435 -75
rect 2395 -205 2435 -195
rect 2505 -75 2545 -65
rect 2505 -195 2515 -75
rect 2535 -195 2545 -75
rect 2505 -205 2545 -195
rect 1815 -285 1835 -205
rect 2225 -220 2245 -205
rect 2225 -230 2265 -220
rect 2225 -250 2235 -230
rect 2255 -250 2265 -230
rect 2225 -260 2265 -250
rect 2395 -285 2415 -205
rect 405 -305 665 -285
rect 955 -305 2415 -285
rect 780 -335 820 -325
rect 185 -360 625 -340
rect -35 -380 -15 -365
rect 185 -380 205 -360
rect 395 -380 415 -360
rect 605 -380 625 -360
rect 780 -355 790 -335
rect 810 -345 820 -335
rect 810 -355 845 -345
rect 780 -365 845 -355
rect 825 -380 845 -365
rect 955 -380 975 -305
rect -55 -390 -15 -380
rect -55 -510 -45 -390
rect -25 -510 -15 -390
rect -55 -520 -15 -510
rect 55 -390 95 -380
rect 55 -510 65 -390
rect 85 -510 95 -390
rect 55 -520 95 -510
rect 165 -390 205 -380
rect 165 -510 175 -390
rect 195 -510 205 -390
rect 165 -520 205 -510
rect 275 -390 315 -380
rect 275 -510 285 -390
rect 305 -510 315 -390
rect 275 -520 315 -510
rect 385 -390 425 -380
rect 385 -510 395 -390
rect 415 -510 425 -390
rect 385 -520 425 -510
rect 495 -390 535 -380
rect 495 -510 505 -390
rect 525 -510 535 -390
rect 495 -520 535 -510
rect 605 -390 645 -380
rect 605 -510 615 -390
rect 635 -510 645 -390
rect 605 -520 645 -510
rect 715 -390 755 -380
rect 715 -510 725 -390
rect 745 -510 755 -390
rect 715 -520 755 -510
rect 825 -390 865 -380
rect 825 -510 835 -390
rect 855 -510 865 -390
rect 825 -520 865 -510
rect 935 -390 975 -380
rect 935 -510 945 -390
rect 965 -510 975 -390
rect 935 -520 975 -510
rect 1045 -335 1085 -325
rect 1045 -355 1055 -335
rect 1075 -355 1085 -335
rect 1045 -390 1085 -355
rect 1045 -510 1055 -390
rect 1075 -510 1085 -390
rect 1045 -520 1085 -510
rect 1155 -380 1175 -305
rect 1395 -335 1475 -325
rect 1395 -355 1405 -335
rect 1465 -355 1475 -335
rect 1395 -365 1475 -355
rect 1395 -380 1415 -365
rect 1595 -380 1615 -305
rect 2565 -325 2585 465
rect 1660 -335 1700 -325
rect 1660 -355 1670 -335
rect 1690 -345 1700 -335
rect 1840 -335 2585 -325
rect 1690 -355 1725 -345
rect 1660 -365 1725 -355
rect 1840 -355 1850 -335
rect 2420 -345 2585 -335
rect 2420 -355 2430 -345
rect 1840 -365 2430 -355
rect 1705 -380 1725 -365
rect 2450 -375 2585 -365
rect 1155 -390 1195 -380
rect 1155 -510 1165 -390
rect 1185 -510 1195 -390
rect 1155 -520 1195 -510
rect 1265 -390 1305 -380
rect 1265 -510 1275 -390
rect 1295 -510 1305 -390
rect 1265 -520 1305 -510
rect 1375 -390 1415 -380
rect 1375 -510 1385 -390
rect 1405 -510 1415 -390
rect 1375 -520 1415 -510
rect 1485 -390 1525 -380
rect 1485 -510 1495 -390
rect 1515 -510 1525 -390
rect 1485 -520 1525 -510
rect 1595 -390 1635 -380
rect 1595 -510 1605 -390
rect 1625 -510 1635 -390
rect 1595 -520 1635 -510
rect 1705 -390 1795 -380
rect 1705 -510 1715 -390
rect 1735 -510 1765 -390
rect 1785 -510 1795 -390
rect 1840 -400 2430 -390
rect 1840 -420 1850 -400
rect 2420 -420 2430 -400
rect 2450 -395 2460 -375
rect 2480 -385 2585 -375
rect 2480 -395 2490 -385
rect 2450 -405 2490 -395
rect 1840 -430 2430 -420
rect 1705 -520 1795 -510
<< viali >>
rect -45 475 -25 595
rect 65 475 85 520
rect 285 475 305 520
rect 505 475 525 520
rect 725 475 745 520
rect 835 475 855 595
rect 1275 475 1295 595
rect 1495 475 1515 595
rect 1490 415 1550 435
rect 1355 335 1375 355
rect -45 175 -25 295
rect 285 175 305 295
rect 505 175 525 295
rect 835 175 855 295
rect 885 175 905 295
rect 935 175 955 295
rect 85 120 145 140
rect 665 120 725 140
rect 985 120 1045 140
rect 1130 45 1190 65
rect 1485 120 1505 140
rect 1715 475 1735 595
rect 1765 475 1785 595
rect 1885 540 2455 560
rect 1885 410 2455 430
rect 1760 375 1800 395
rect 1800 375 1820 395
rect 1595 175 1615 295
rect 1695 175 1715 295
rect 2105 250 2125 295
rect 2215 250 2235 295
rect 2515 175 2535 295
rect 1290 10 1330 30
rect 1330 10 1350 30
rect 1420 10 1440 30
rect 1525 20 1585 40
rect -45 -195 -25 -75
rect 285 -195 305 -75
rect 505 -195 525 -75
rect 835 -195 855 -75
rect 885 -195 905 -75
rect 935 -195 955 -75
rect 1265 -120 1285 -75
rect 1595 -195 1615 -75
rect 195 -255 255 -235
rect 555 -255 615 -235
rect 1695 -195 1715 -75
rect 2105 -195 2125 -150
rect 2515 -195 2535 -75
rect -45 -510 -25 -390
rect 65 -435 85 -390
rect 285 -435 305 -390
rect 505 -435 525 -390
rect 725 -435 745 -390
rect 835 -510 855 -390
rect 1405 -355 1465 -335
rect 1275 -510 1295 -390
rect 1495 -510 1515 -390
rect 1715 -510 1735 -390
rect 1850 -420 2420 -400
<< metal1 >>
rect -60 595 1795 605
rect -60 475 -45 595
rect -25 545 835 595
rect -25 475 -15 545
rect -60 465 -15 475
rect 55 520 755 530
rect 55 475 65 520
rect 85 475 285 520
rect 305 475 505 520
rect 525 475 720 520
rect 750 475 755 520
rect 55 465 755 475
rect 825 475 835 545
rect 855 475 1275 595
rect 1295 475 1495 595
rect 1515 475 1715 595
rect 1735 475 1765 595
rect 1785 570 1795 595
rect 1785 560 2465 570
rect 1785 540 1885 560
rect 2455 540 2465 560
rect 1785 475 2465 540
rect 825 465 2465 475
rect 1480 435 1560 445
rect 1480 415 1490 435
rect 1550 425 1560 435
rect 1875 440 2465 465
rect 1875 430 2545 440
rect 1550 415 1705 425
rect 1480 405 1705 415
rect 1875 410 1885 430
rect 2455 410 2545 430
rect 1345 355 1385 365
rect 1345 335 1355 355
rect 1375 345 1385 355
rect 1685 345 1705 405
rect 1750 395 1830 405
rect 1875 400 2545 410
rect 1750 375 1760 395
rect 1820 385 1830 395
rect 1820 375 2245 385
rect 1750 360 2245 375
rect 1375 335 1665 345
rect 1345 325 1665 335
rect 1685 325 2135 345
rect -80 295 1630 305
rect -80 175 -45 295
rect -25 220 285 295
rect -25 175 60 220
rect 90 175 285 220
rect 305 175 505 295
rect 525 175 835 295
rect 855 175 885 295
rect 905 175 935 295
rect 955 175 1595 295
rect 1615 175 1630 295
rect -80 165 1630 175
rect 75 140 735 150
rect 75 120 85 140
rect 145 120 665 140
rect 725 120 735 140
rect 75 110 735 120
rect 975 140 1540 150
rect 975 120 985 140
rect 1045 130 1485 140
rect 1045 120 1055 130
rect 975 110 1055 120
rect 1475 120 1485 130
rect 1505 120 1540 140
rect 1475 110 1540 120
rect 1120 65 1200 75
rect 1120 55 1130 65
rect -80 45 1130 55
rect 1190 45 1200 65
rect -80 35 1200 45
rect 1515 50 1540 110
rect 1515 40 1595 50
rect 1280 30 1360 40
rect 1280 20 1290 30
rect -80 10 1290 20
rect 1350 10 1360 30
rect -80 0 1360 10
rect 1410 30 1450 40
rect 1410 10 1420 30
rect 1440 10 1450 30
rect 1515 20 1525 40
rect 1585 20 1595 40
rect 1515 10 1595 20
rect 1410 0 1450 10
rect 1415 -25 1430 0
rect 1280 -40 1430 -25
rect 1280 -65 1295 -40
rect -80 -75 1185 -65
rect -80 -195 -45 -75
rect -25 -195 285 -75
rect 305 -195 505 -75
rect 525 -120 720 -75
rect 750 -120 835 -75
rect 525 -195 835 -120
rect 855 -195 885 -75
rect 905 -195 935 -75
rect 955 -145 1185 -75
rect 1255 -75 1295 -65
rect 1255 -120 1265 -75
rect 1285 -120 1295 -75
rect 1255 -130 1295 -120
rect 1365 -75 1630 -65
rect 1365 -145 1595 -75
rect 955 -195 1595 -145
rect 1615 -195 1630 -75
rect -80 -205 1630 -195
rect 1645 -220 1665 325
rect 1685 295 2025 305
rect 1685 175 1695 295
rect 1715 215 2025 295
rect 2095 295 2135 325
rect 2095 250 2105 295
rect 2125 250 2135 295
rect 2095 240 2135 250
rect 2205 295 2245 360
rect 2205 250 2215 295
rect 2235 250 2245 295
rect 2205 240 2245 250
rect 2505 295 2545 400
rect 2505 215 2515 295
rect 1715 175 2515 215
rect 2535 175 2545 295
rect 1685 165 2545 175
rect 1685 -75 2545 -65
rect 1685 -195 1695 -75
rect 1715 -115 2515 -75
rect 1715 -195 2025 -115
rect 1685 -205 2025 -195
rect 2095 -150 2135 -140
rect 2095 -195 2105 -150
rect 2125 -195 2135 -150
rect 2095 -220 2135 -195
rect 2205 -195 2515 -115
rect 2535 -195 2545 -75
rect 2205 -205 2545 -195
rect 185 -235 625 -225
rect 185 -255 195 -235
rect 255 -255 555 -235
rect 615 -255 625 -235
rect 185 -265 625 -255
rect 1460 -235 2135 -220
rect 1460 -325 1475 -235
rect 1395 -335 1475 -325
rect 1395 -355 1405 -335
rect 1465 -355 1475 -335
rect 1395 -365 1475 -355
rect -55 -390 -15 -380
rect -55 -510 -45 -390
rect -25 -460 -15 -390
rect 55 -390 755 -380
rect 55 -435 60 -390
rect 90 -435 285 -390
rect 305 -435 505 -390
rect 525 -435 725 -390
rect 745 -435 755 -390
rect 55 -445 755 -435
rect 825 -390 1795 -380
rect 825 -460 835 -390
rect -25 -510 835 -460
rect 855 -510 1275 -390
rect 1295 -510 1495 -390
rect 1515 -510 1715 -390
rect 1735 -400 2430 -390
rect 1735 -420 1850 -400
rect 2420 -420 2430 -400
rect 1735 -430 2430 -420
rect 1735 -510 1795 -430
rect -55 -520 1795 -510
<< via1 >>
rect 720 475 725 520
rect 725 475 745 520
rect 745 475 750 520
rect 60 175 90 220
rect 720 -120 750 -75
rect 60 -435 65 -390
rect 65 -435 85 -390
rect 85 -435 90 -390
<< metal2 >>
rect 715 520 755 530
rect 715 475 720 520
rect 750 475 755 520
rect 55 220 95 230
rect 55 175 60 220
rect 90 175 95 220
rect 55 -390 95 175
rect 715 -75 755 475
rect 715 -120 720 -75
rect 750 -120 755 -75
rect 715 -130 755 -120
rect 55 -435 60 -390
rect 90 -435 95 -390
rect 55 -445 95 -435
<< labels >>
rlabel metal1 -80 235 -80 235 7 VP
port 0 w
rlabel metal1 -80 -135 -80 -135 7 VN
port 1 w
rlabel metal1 -80 45 -80 45 7 V1
port 2 w
rlabel metal1 -80 10 -80 10 7 V2
port 3 w
rlabel locali 2585 80 2585 80 3 Vout
port 4 e
rlabel locali 2585 -375 2585 -375 3 nVout
port 5 e
<< end >>
