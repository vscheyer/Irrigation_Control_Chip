magic
tech sky130A
timestamp 1620340807
<< nwell >>
rect -70 195 345 355
<< nmos >>
rect 0 20 15 120
rect 65 20 80 120
rect 210 20 225 120
<< pmos >>
rect 0 225 15 325
rect 65 225 80 325
rect 210 225 225 325
<< ndiff >>
rect -50 105 0 120
rect -50 35 -35 105
rect -15 35 0 105
rect -50 20 0 35
rect 15 105 65 120
rect 15 35 30 105
rect 50 35 65 105
rect 15 20 65 35
rect 80 105 130 120
rect 80 35 95 105
rect 115 35 130 105
rect 80 20 130 35
rect 160 105 210 120
rect 160 35 175 105
rect 195 35 210 105
rect 160 20 210 35
rect 225 105 275 120
rect 225 35 240 105
rect 260 35 275 105
rect 225 20 275 35
<< pdiff >>
rect -50 310 0 325
rect -50 240 -35 310
rect -15 240 0 310
rect -50 225 0 240
rect 15 310 65 325
rect 15 240 30 310
rect 50 240 65 310
rect 15 225 65 240
rect 80 310 130 325
rect 80 240 95 310
rect 115 240 130 310
rect 80 225 130 240
rect 160 310 210 325
rect 160 240 175 310
rect 195 240 210 310
rect 160 225 210 240
rect 225 310 275 325
rect 225 240 240 310
rect 260 240 275 310
rect 225 225 275 240
<< ndiffc >>
rect -35 35 -15 105
rect 30 35 50 105
rect 95 35 115 105
rect 175 35 195 105
rect 240 35 260 105
<< pdiffc >>
rect -35 240 -15 310
rect 30 240 50 310
rect 95 240 115 310
rect 175 240 195 310
rect 240 240 260 310
<< psubdiff >>
rect 275 105 325 120
rect 275 35 290 105
rect 310 35 325 105
rect 275 20 325 35
<< nsubdiff >>
rect 275 310 325 325
rect 275 240 290 310
rect 310 240 325 310
rect 275 225 325 240
<< psubdiffcont >>
rect 290 35 310 105
<< nsubdiffcont >>
rect 290 240 310 310
<< poly >>
rect -25 370 15 380
rect -25 350 -15 370
rect 5 350 15 370
rect -25 340 15 350
rect 0 325 15 340
rect 65 325 80 340
rect 210 325 225 340
rect 0 210 15 225
rect 65 215 80 225
rect 210 215 225 225
rect 65 200 225 215
rect 65 185 80 200
rect 0 170 80 185
rect 210 175 225 200
rect 0 120 15 170
rect 145 160 185 170
rect 145 145 155 160
rect 65 140 155 145
rect 175 140 185 160
rect 65 130 185 140
rect 210 165 250 175
rect 210 145 220 165
rect 240 145 250 165
rect 210 135 250 145
rect 65 120 80 130
rect 210 120 225 135
rect 0 5 15 20
rect 65 5 80 20
rect 210 5 225 20
<< polycont >>
rect -15 350 5 370
rect 155 140 175 160
rect 220 145 240 165
<< locali >>
rect -25 370 15 380
rect -25 350 -15 370
rect 5 360 15 370
rect 5 350 185 360
rect -25 340 185 350
rect 165 320 185 340
rect -45 310 -5 320
rect -45 240 -35 310
rect -15 240 -5 310
rect -45 230 -5 240
rect 20 310 60 320
rect 20 240 30 310
rect 50 240 60 310
rect 20 230 60 240
rect 85 310 125 320
rect 85 240 95 310
rect 115 240 125 310
rect 85 230 125 240
rect 165 310 205 320
rect 165 240 175 310
rect 195 240 205 310
rect 165 230 205 240
rect 230 310 345 320
rect 230 240 240 310
rect 260 240 290 310
rect 310 240 345 310
rect 230 230 345 240
rect -45 115 -25 230
rect 20 115 40 230
rect 85 115 105 230
rect 165 170 185 230
rect 145 160 185 170
rect 145 140 155 160
rect 175 140 185 160
rect 145 130 185 140
rect 210 165 250 175
rect 210 145 220 165
rect 240 155 250 165
rect 240 145 345 155
rect 210 135 345 145
rect 165 115 185 130
rect -45 105 -5 115
rect -45 35 -35 105
rect -15 35 -5 105
rect -45 25 -5 35
rect 20 105 60 115
rect 20 35 30 105
rect 50 35 60 105
rect 20 25 60 35
rect 85 105 125 115
rect 85 35 95 105
rect 115 35 125 105
rect 85 25 125 35
rect 165 105 205 115
rect 165 35 175 105
rect 195 35 205 105
rect 165 25 205 35
rect 230 105 345 115
rect 230 35 240 105
rect 260 35 290 105
rect 310 35 345 105
rect 230 25 345 35
rect -45 5 -25 25
rect 20 5 40 25
rect 85 5 105 25
<< labels >>
rlabel locali 345 275 345 275 3 VP
port 0 e
rlabel locali 345 70 345 70 3 VN
port 1 e
rlabel locali 95 5 95 5 5 A
port 2 s
rlabel locali -35 5 -35 5 5 B
port 3 s
rlabel locali 345 145 345 145 3 C
port 4 e
rlabel locali 30 5 30 5 5 Out
port 5 s
<< end >>
