magic
tech sky130A
magscale 1 2
timestamp 1620791022
<< locali >>
rect 13185 2839 13219 3077
<< viali >>
rect 27261 29733 27295 29767
rect 1409 29665 1443 29699
rect 9597 29665 9631 29699
rect 19349 29665 19383 29699
rect 1593 29461 1627 29495
rect 9781 29461 9815 29495
rect 27169 29461 27203 29495
rect 27997 17017 28031 17051
rect 28181 17017 28215 17051
rect 14933 15521 14967 15555
rect 14841 15317 14875 15351
rect 1409 14909 1443 14943
rect 12357 14909 12391 14943
rect 12817 14909 12851 14943
rect 13001 14909 13035 14943
rect 13093 14909 13127 14943
rect 13185 14909 13219 14943
rect 1593 14773 1627 14807
rect 12265 14773 12299 14807
rect 13461 14773 13495 14807
rect 12173 14433 12207 14467
rect 12633 14433 12667 14467
rect 12817 14433 12851 14467
rect 12909 14433 12943 14467
rect 13001 14433 13035 14467
rect 12081 14365 12115 14399
rect 13277 14229 13311 14263
rect 11069 13889 11103 13923
rect 10977 13821 11011 13855
rect 11161 13821 11195 13855
rect 13194 13821 13228 13855
rect 13461 13821 13495 13855
rect 13921 13821 13955 13855
rect 14188 13753 14222 13787
rect 12081 13685 12115 13719
rect 15301 13685 15335 13719
rect 11713 13481 11747 13515
rect 10793 13345 10827 13379
rect 10885 13345 10919 13379
rect 11989 13345 12023 13379
rect 12173 13345 12207 13379
rect 13277 13345 13311 13379
rect 13461 13345 13495 13379
rect 11897 13277 11931 13311
rect 12081 13277 12115 13311
rect 13185 13277 13219 13311
rect 13645 13141 13679 13175
rect 13553 12937 13587 12971
rect 14381 12937 14415 12971
rect 10977 12733 11011 12767
rect 12173 12733 12207 12767
rect 14013 12733 14047 12767
rect 12440 12665 12474 12699
rect 14197 12665 14231 12699
rect 11069 12597 11103 12631
rect 12633 12393 12667 12427
rect 10508 12257 10542 12291
rect 12817 12257 12851 12291
rect 13093 12257 13127 12291
rect 13645 12257 13679 12291
rect 14749 12257 14783 12291
rect 14933 12257 14967 12291
rect 10241 12189 10275 12223
rect 12909 12189 12943 12223
rect 13001 12189 13035 12223
rect 11621 12053 11655 12087
rect 13829 12053 13863 12087
rect 14933 12053 14967 12087
rect 12817 11849 12851 11883
rect 13277 11849 13311 11883
rect 13645 11849 13679 11883
rect 9781 11781 9815 11815
rect 12357 11713 12391 11747
rect 14933 11713 14967 11747
rect 9873 11645 9907 11679
rect 10333 11645 10367 11679
rect 10517 11645 10551 11679
rect 12081 11645 12115 11679
rect 12265 11645 12299 11679
rect 12449 11645 12483 11679
rect 12633 11645 12667 11679
rect 13461 11645 13495 11679
rect 13645 11645 13679 11679
rect 14657 11645 14691 11679
rect 15669 11645 15703 11679
rect 10701 11509 10735 11543
rect 14289 11509 14323 11543
rect 14749 11509 14783 11543
rect 15577 11509 15611 11543
rect 11529 11305 11563 11339
rect 12725 11305 12759 11339
rect 13553 11305 13587 11339
rect 16129 11305 16163 11339
rect 10802 11237 10836 11271
rect 12541 11237 12575 11271
rect 14994 11237 15028 11271
rect 11069 11169 11103 11203
rect 11713 11169 11747 11203
rect 11897 11169 11931 11203
rect 12357 11169 12391 11203
rect 13645 11169 13679 11203
rect 13829 11169 13863 11203
rect 14749 11169 14783 11203
rect 9689 10965 9723 10999
rect 13369 10965 13403 10999
rect 9965 10761 9999 10795
rect 10977 10761 11011 10795
rect 11161 10761 11195 10795
rect 12357 10761 12391 10795
rect 12541 10761 12575 10795
rect 12817 10761 12851 10795
rect 13461 10761 13495 10795
rect 14289 10761 14323 10795
rect 15761 10761 15795 10795
rect 15945 10761 15979 10795
rect 12449 10693 12483 10727
rect 15301 10625 15335 10659
rect 10149 10557 10183 10591
rect 12081 10557 12115 10591
rect 13277 10557 13311 10591
rect 13461 10557 13495 10591
rect 13921 10557 13955 10591
rect 14289 10557 14323 10591
rect 15117 10557 15151 10591
rect 10333 10489 10367 10523
rect 10793 10489 10827 10523
rect 16129 10489 16163 10523
rect 10998 10421 11032 10455
rect 12173 10421 12207 10455
rect 14105 10421 14139 10455
rect 14933 10421 14967 10455
rect 15924 10421 15958 10455
rect 13093 10217 13127 10251
rect 16129 10217 16163 10251
rect 12725 10149 12759 10183
rect 10313 10081 10347 10115
rect 12081 10081 12115 10115
rect 12265 10081 12299 10115
rect 12909 10081 12943 10115
rect 13645 10081 13679 10115
rect 15005 10081 15039 10115
rect 10057 10013 10091 10047
rect 14749 10013 14783 10047
rect 13829 9945 13863 9979
rect 11437 9877 11471 9911
rect 11897 9877 11931 9911
rect 12173 9673 12207 9707
rect 13921 9673 13955 9707
rect 9781 9537 9815 9571
rect 12081 9537 12115 9571
rect 14473 9537 14507 9571
rect 15301 9537 15335 9571
rect 12265 9469 12299 9503
rect 12357 9469 12391 9503
rect 13829 9469 13863 9503
rect 14013 9469 14047 9503
rect 15485 9469 15519 9503
rect 15577 9469 15611 9503
rect 16037 9469 16071 9503
rect 10048 9401 10082 9435
rect 14657 9401 14691 9435
rect 14841 9401 14875 9435
rect 15301 9401 15335 9435
rect 11161 9333 11195 9367
rect 16129 9333 16163 9367
rect 10425 9129 10459 9163
rect 10977 9129 11011 9163
rect 11161 9129 11195 9163
rect 15016 9061 15050 9095
rect 10517 8993 10551 9027
rect 11158 8993 11192 9027
rect 11621 8993 11655 9027
rect 12081 8993 12115 9027
rect 14749 8993 14783 9027
rect 13369 8857 13403 8891
rect 11529 8789 11563 8823
rect 16129 8789 16163 8823
rect 10885 8585 10919 8619
rect 12173 8585 12207 8619
rect 15301 8449 15335 8483
rect 10977 8381 11011 8415
rect 12081 8381 12115 8415
rect 12265 8381 12299 8415
rect 13737 8381 13771 8415
rect 13829 8381 13863 8415
rect 14565 8381 14599 8415
rect 14657 8381 14691 8415
rect 15209 8381 15243 8415
rect 15393 8381 15427 8415
rect 13277 8041 13311 8075
rect 12633 7973 12667 8007
rect 14994 7973 15028 8007
rect 10793 7905 10827 7939
rect 11897 7905 11931 7939
rect 12541 7905 12575 7939
rect 12817 7905 12851 7939
rect 13461 7905 13495 7939
rect 10609 7837 10643 7871
rect 11713 7837 11747 7871
rect 14749 7837 14783 7871
rect 10977 7701 11011 7735
rect 12081 7701 12115 7735
rect 12541 7701 12575 7735
rect 16129 7701 16163 7735
rect 9781 7497 9815 7531
rect 12265 7497 12299 7531
rect 14749 7497 14783 7531
rect 10894 7293 10928 7327
rect 11161 7293 11195 7327
rect 14105 7293 14139 7327
rect 14289 7293 14323 7327
rect 14381 7293 14415 7327
rect 14473 7293 14507 7327
rect 15209 7293 15243 7327
rect 15393 7293 15427 7327
rect 12081 7225 12115 7259
rect 12297 7225 12331 7259
rect 13553 7225 13587 7259
rect 15301 7225 15335 7259
rect 12449 7157 12483 7191
rect 13461 7157 13495 7191
rect 11468 6885 11502 6919
rect 11713 6817 11747 6851
rect 12265 6817 12299 6851
rect 12449 6817 12483 6851
rect 12817 6817 12851 6851
rect 13461 6817 13495 6851
rect 13645 6817 13679 6851
rect 14933 6817 14967 6851
rect 15393 6817 15427 6851
rect 15577 6817 15611 6851
rect 12541 6749 12575 6783
rect 12633 6749 12667 6783
rect 13001 6681 13035 6715
rect 10333 6613 10367 6647
rect 13737 6613 13771 6647
rect 14749 6613 14783 6647
rect 15393 6613 15427 6647
rect 11161 6409 11195 6443
rect 12081 6409 12115 6443
rect 13277 6409 13311 6443
rect 10149 6205 10183 6239
rect 10793 6205 10827 6239
rect 12219 6205 12253 6239
rect 12632 6205 12666 6239
rect 12725 6205 12759 6239
rect 13369 6205 13403 6239
rect 13829 6205 13863 6239
rect 14096 6205 14130 6239
rect 10977 6137 11011 6171
rect 12357 6137 12391 6171
rect 12449 6137 12483 6171
rect 10333 6069 10367 6103
rect 15209 6069 15243 6103
rect 11069 5865 11103 5899
rect 14841 5865 14875 5899
rect 10885 5797 10919 5831
rect 11529 5797 11563 5831
rect 11713 5797 11747 5831
rect 10701 5729 10735 5763
rect 11897 5729 11931 5763
rect 12541 5729 12575 5763
rect 12725 5729 12759 5763
rect 13277 5729 13311 5763
rect 13461 5729 13495 5763
rect 14933 5729 14967 5763
rect 12357 5661 12391 5695
rect 13645 5661 13679 5695
rect 12265 5321 12299 5355
rect 13277 5321 13311 5355
rect 12541 5185 12575 5219
rect 11161 5117 11195 5151
rect 12449 5117 12483 5151
rect 12633 5117 12667 5151
rect 12725 5117 12759 5151
rect 13461 5117 13495 5151
rect 13553 5117 13587 5151
rect 13737 5117 13771 5151
rect 13829 5117 13863 5151
rect 14289 5117 14323 5151
rect 14473 5117 14507 5151
rect 15945 5117 15979 5151
rect 14381 5049 14415 5083
rect 11069 4981 11103 5015
rect 15853 4981 15887 5015
rect 11897 4777 11931 4811
rect 12718 4777 12752 4811
rect 13553 4777 13587 4811
rect 13829 4777 13863 4811
rect 16221 4777 16255 4811
rect 10784 4709 10818 4743
rect 12817 4709 12851 4743
rect 13645 4709 13679 4743
rect 10057 4641 10091 4675
rect 10517 4641 10551 4675
rect 12541 4641 12575 4675
rect 12633 4641 12667 4675
rect 13461 4641 13495 4675
rect 14749 4641 14783 4675
rect 16313 4641 16347 4675
rect 16405 4573 16439 4607
rect 13277 4505 13311 4539
rect 9965 4437 9999 4471
rect 14841 4437 14875 4471
rect 15853 4437 15887 4471
rect 14381 4233 14415 4267
rect 16405 4233 16439 4267
rect 12399 4097 12433 4131
rect 10977 4029 11011 4063
rect 11161 4029 11195 4063
rect 12173 4029 12207 4063
rect 12541 4029 12575 4063
rect 13001 4029 13035 4063
rect 15025 4029 15059 4063
rect 15292 4029 15326 4063
rect 13246 3961 13280 3995
rect 11069 3893 11103 3927
rect 12265 3893 12299 3927
rect 12449 3893 12483 3927
rect 12449 3689 12483 3723
rect 15117 3689 15151 3723
rect 15485 3689 15519 3723
rect 10854 3621 10888 3655
rect 10609 3553 10643 3587
rect 13562 3553 13596 3587
rect 13829 3553 13863 3587
rect 15577 3553 15611 3587
rect 15669 3485 15703 3519
rect 11989 3349 12023 3383
rect 12357 3145 12391 3179
rect 19901 3145 19935 3179
rect 27905 3145 27939 3179
rect 13185 3077 13219 3111
rect 13921 3077 13955 3111
rect 12173 2941 12207 2975
rect 12357 2941 12391 2975
rect 12725 2941 12759 2975
rect 13461 2941 13495 2975
rect 14105 2941 14139 2975
rect 19993 2941 20027 2975
rect 27813 2941 27847 2975
rect 12633 2805 12667 2839
rect 13185 2805 13219 2839
rect 13277 2805 13311 2839
rect 1593 2601 1627 2635
rect 20729 2601 20763 2635
rect 27353 2601 27387 2635
rect 1409 2465 1443 2499
rect 20913 2465 20947 2499
rect 27169 2465 27203 2499
<< metal1 >>
rect 1104 29946 28888 29968
rect 1104 29894 10243 29946
rect 10295 29894 10307 29946
rect 10359 29894 10371 29946
rect 10423 29894 10435 29946
rect 10487 29894 19504 29946
rect 19556 29894 19568 29946
rect 19620 29894 19632 29946
rect 19684 29894 19696 29946
rect 19748 29894 28888 29946
rect 1104 29872 28888 29894
rect 27249 29767 27307 29773
rect 27249 29733 27261 29767
rect 27295 29764 27307 29767
rect 29454 29764 29460 29776
rect 27295 29736 29460 29764
rect 27295 29733 27307 29736
rect 27249 29727 27307 29733
rect 29454 29724 29460 29736
rect 29512 29724 29518 29776
rect 1394 29696 1400 29708
rect 1355 29668 1400 29696
rect 1394 29656 1400 29668
rect 1452 29656 1458 29708
rect 9214 29656 9220 29708
rect 9272 29696 9278 29708
rect 9585 29699 9643 29705
rect 9585 29696 9597 29699
rect 9272 29668 9597 29696
rect 9272 29656 9278 29668
rect 9585 29665 9597 29668
rect 9631 29665 9643 29699
rect 19334 29696 19340 29708
rect 19295 29668 19340 29696
rect 9585 29659 9643 29665
rect 19334 29656 19340 29668
rect 19392 29656 19398 29708
rect 1578 29492 1584 29504
rect 1539 29464 1584 29492
rect 1578 29452 1584 29464
rect 1636 29452 1642 29504
rect 9766 29492 9772 29504
rect 9727 29464 9772 29492
rect 9766 29452 9772 29464
rect 9824 29452 9830 29504
rect 14734 29452 14740 29504
rect 14792 29492 14798 29504
rect 27157 29495 27215 29501
rect 27157 29492 27169 29495
rect 14792 29464 27169 29492
rect 14792 29452 14798 29464
rect 27157 29461 27169 29464
rect 27203 29461 27215 29495
rect 27157 29455 27215 29461
rect 1104 29402 28888 29424
rect 1104 29350 5612 29402
rect 5664 29350 5676 29402
rect 5728 29350 5740 29402
rect 5792 29350 5804 29402
rect 5856 29350 14874 29402
rect 14926 29350 14938 29402
rect 14990 29350 15002 29402
rect 15054 29350 15066 29402
rect 15118 29350 24135 29402
rect 24187 29350 24199 29402
rect 24251 29350 24263 29402
rect 24315 29350 24327 29402
rect 24379 29350 28888 29402
rect 1104 29328 28888 29350
rect 1104 28858 28888 28880
rect 1104 28806 10243 28858
rect 10295 28806 10307 28858
rect 10359 28806 10371 28858
rect 10423 28806 10435 28858
rect 10487 28806 19504 28858
rect 19556 28806 19568 28858
rect 19620 28806 19632 28858
rect 19684 28806 19696 28858
rect 19748 28806 28888 28858
rect 1104 28784 28888 28806
rect 1104 28314 28888 28336
rect 1104 28262 5612 28314
rect 5664 28262 5676 28314
rect 5728 28262 5740 28314
rect 5792 28262 5804 28314
rect 5856 28262 14874 28314
rect 14926 28262 14938 28314
rect 14990 28262 15002 28314
rect 15054 28262 15066 28314
rect 15118 28262 24135 28314
rect 24187 28262 24199 28314
rect 24251 28262 24263 28314
rect 24315 28262 24327 28314
rect 24379 28262 28888 28314
rect 1104 28240 28888 28262
rect 1104 27770 28888 27792
rect 1104 27718 10243 27770
rect 10295 27718 10307 27770
rect 10359 27718 10371 27770
rect 10423 27718 10435 27770
rect 10487 27718 19504 27770
rect 19556 27718 19568 27770
rect 19620 27718 19632 27770
rect 19684 27718 19696 27770
rect 19748 27718 28888 27770
rect 1104 27696 28888 27718
rect 1104 27226 28888 27248
rect 1104 27174 5612 27226
rect 5664 27174 5676 27226
rect 5728 27174 5740 27226
rect 5792 27174 5804 27226
rect 5856 27174 14874 27226
rect 14926 27174 14938 27226
rect 14990 27174 15002 27226
rect 15054 27174 15066 27226
rect 15118 27174 24135 27226
rect 24187 27174 24199 27226
rect 24251 27174 24263 27226
rect 24315 27174 24327 27226
rect 24379 27174 28888 27226
rect 1104 27152 28888 27174
rect 1104 26682 28888 26704
rect 1104 26630 10243 26682
rect 10295 26630 10307 26682
rect 10359 26630 10371 26682
rect 10423 26630 10435 26682
rect 10487 26630 19504 26682
rect 19556 26630 19568 26682
rect 19620 26630 19632 26682
rect 19684 26630 19696 26682
rect 19748 26630 28888 26682
rect 1104 26608 28888 26630
rect 1104 26138 28888 26160
rect 1104 26086 5612 26138
rect 5664 26086 5676 26138
rect 5728 26086 5740 26138
rect 5792 26086 5804 26138
rect 5856 26086 14874 26138
rect 14926 26086 14938 26138
rect 14990 26086 15002 26138
rect 15054 26086 15066 26138
rect 15118 26086 24135 26138
rect 24187 26086 24199 26138
rect 24251 26086 24263 26138
rect 24315 26086 24327 26138
rect 24379 26086 28888 26138
rect 1104 26064 28888 26086
rect 1104 25594 28888 25616
rect 1104 25542 10243 25594
rect 10295 25542 10307 25594
rect 10359 25542 10371 25594
rect 10423 25542 10435 25594
rect 10487 25542 19504 25594
rect 19556 25542 19568 25594
rect 19620 25542 19632 25594
rect 19684 25542 19696 25594
rect 19748 25542 28888 25594
rect 1104 25520 28888 25542
rect 1104 25050 28888 25072
rect 1104 24998 5612 25050
rect 5664 24998 5676 25050
rect 5728 24998 5740 25050
rect 5792 24998 5804 25050
rect 5856 24998 14874 25050
rect 14926 24998 14938 25050
rect 14990 24998 15002 25050
rect 15054 24998 15066 25050
rect 15118 24998 24135 25050
rect 24187 24998 24199 25050
rect 24251 24998 24263 25050
rect 24315 24998 24327 25050
rect 24379 24998 28888 25050
rect 1104 24976 28888 24998
rect 1104 24506 28888 24528
rect 1104 24454 10243 24506
rect 10295 24454 10307 24506
rect 10359 24454 10371 24506
rect 10423 24454 10435 24506
rect 10487 24454 19504 24506
rect 19556 24454 19568 24506
rect 19620 24454 19632 24506
rect 19684 24454 19696 24506
rect 19748 24454 28888 24506
rect 1104 24432 28888 24454
rect 1104 23962 28888 23984
rect 1104 23910 5612 23962
rect 5664 23910 5676 23962
rect 5728 23910 5740 23962
rect 5792 23910 5804 23962
rect 5856 23910 14874 23962
rect 14926 23910 14938 23962
rect 14990 23910 15002 23962
rect 15054 23910 15066 23962
rect 15118 23910 24135 23962
rect 24187 23910 24199 23962
rect 24251 23910 24263 23962
rect 24315 23910 24327 23962
rect 24379 23910 28888 23962
rect 1104 23888 28888 23910
rect 1104 23418 28888 23440
rect 1104 23366 10243 23418
rect 10295 23366 10307 23418
rect 10359 23366 10371 23418
rect 10423 23366 10435 23418
rect 10487 23366 19504 23418
rect 19556 23366 19568 23418
rect 19620 23366 19632 23418
rect 19684 23366 19696 23418
rect 19748 23366 28888 23418
rect 1104 23344 28888 23366
rect 1104 22874 28888 22896
rect 1104 22822 5612 22874
rect 5664 22822 5676 22874
rect 5728 22822 5740 22874
rect 5792 22822 5804 22874
rect 5856 22822 14874 22874
rect 14926 22822 14938 22874
rect 14990 22822 15002 22874
rect 15054 22822 15066 22874
rect 15118 22822 24135 22874
rect 24187 22822 24199 22874
rect 24251 22822 24263 22874
rect 24315 22822 24327 22874
rect 24379 22822 28888 22874
rect 1104 22800 28888 22822
rect 1104 22330 28888 22352
rect 1104 22278 10243 22330
rect 10295 22278 10307 22330
rect 10359 22278 10371 22330
rect 10423 22278 10435 22330
rect 10487 22278 19504 22330
rect 19556 22278 19568 22330
rect 19620 22278 19632 22330
rect 19684 22278 19696 22330
rect 19748 22278 28888 22330
rect 1104 22256 28888 22278
rect 1104 21786 28888 21808
rect 1104 21734 5612 21786
rect 5664 21734 5676 21786
rect 5728 21734 5740 21786
rect 5792 21734 5804 21786
rect 5856 21734 14874 21786
rect 14926 21734 14938 21786
rect 14990 21734 15002 21786
rect 15054 21734 15066 21786
rect 15118 21734 24135 21786
rect 24187 21734 24199 21786
rect 24251 21734 24263 21786
rect 24315 21734 24327 21786
rect 24379 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 10243 21242
rect 10295 21190 10307 21242
rect 10359 21190 10371 21242
rect 10423 21190 10435 21242
rect 10487 21190 19504 21242
rect 19556 21190 19568 21242
rect 19620 21190 19632 21242
rect 19684 21190 19696 21242
rect 19748 21190 28888 21242
rect 1104 21168 28888 21190
rect 1104 20698 28888 20720
rect 1104 20646 5612 20698
rect 5664 20646 5676 20698
rect 5728 20646 5740 20698
rect 5792 20646 5804 20698
rect 5856 20646 14874 20698
rect 14926 20646 14938 20698
rect 14990 20646 15002 20698
rect 15054 20646 15066 20698
rect 15118 20646 24135 20698
rect 24187 20646 24199 20698
rect 24251 20646 24263 20698
rect 24315 20646 24327 20698
rect 24379 20646 28888 20698
rect 1104 20624 28888 20646
rect 1104 20154 28888 20176
rect 1104 20102 10243 20154
rect 10295 20102 10307 20154
rect 10359 20102 10371 20154
rect 10423 20102 10435 20154
rect 10487 20102 19504 20154
rect 19556 20102 19568 20154
rect 19620 20102 19632 20154
rect 19684 20102 19696 20154
rect 19748 20102 28888 20154
rect 1104 20080 28888 20102
rect 1104 19610 28888 19632
rect 1104 19558 5612 19610
rect 5664 19558 5676 19610
rect 5728 19558 5740 19610
rect 5792 19558 5804 19610
rect 5856 19558 14874 19610
rect 14926 19558 14938 19610
rect 14990 19558 15002 19610
rect 15054 19558 15066 19610
rect 15118 19558 24135 19610
rect 24187 19558 24199 19610
rect 24251 19558 24263 19610
rect 24315 19558 24327 19610
rect 24379 19558 28888 19610
rect 1104 19536 28888 19558
rect 1104 19066 28888 19088
rect 1104 19014 10243 19066
rect 10295 19014 10307 19066
rect 10359 19014 10371 19066
rect 10423 19014 10435 19066
rect 10487 19014 19504 19066
rect 19556 19014 19568 19066
rect 19620 19014 19632 19066
rect 19684 19014 19696 19066
rect 19748 19014 28888 19066
rect 1104 18992 28888 19014
rect 1104 18522 28888 18544
rect 1104 18470 5612 18522
rect 5664 18470 5676 18522
rect 5728 18470 5740 18522
rect 5792 18470 5804 18522
rect 5856 18470 14874 18522
rect 14926 18470 14938 18522
rect 14990 18470 15002 18522
rect 15054 18470 15066 18522
rect 15118 18470 24135 18522
rect 24187 18470 24199 18522
rect 24251 18470 24263 18522
rect 24315 18470 24327 18522
rect 24379 18470 28888 18522
rect 1104 18448 28888 18470
rect 1104 17978 28888 18000
rect 1104 17926 10243 17978
rect 10295 17926 10307 17978
rect 10359 17926 10371 17978
rect 10423 17926 10435 17978
rect 10487 17926 19504 17978
rect 19556 17926 19568 17978
rect 19620 17926 19632 17978
rect 19684 17926 19696 17978
rect 19748 17926 28888 17978
rect 1104 17904 28888 17926
rect 1104 17434 28888 17456
rect 1104 17382 5612 17434
rect 5664 17382 5676 17434
rect 5728 17382 5740 17434
rect 5792 17382 5804 17434
rect 5856 17382 14874 17434
rect 14926 17382 14938 17434
rect 14990 17382 15002 17434
rect 15054 17382 15066 17434
rect 15118 17382 24135 17434
rect 24187 17382 24199 17434
rect 24251 17382 24263 17434
rect 24315 17382 24327 17434
rect 24379 17382 28888 17434
rect 1104 17360 28888 17382
rect 27982 17048 27988 17060
rect 27943 17020 27988 17048
rect 27982 17008 27988 17020
rect 28040 17008 28046 17060
rect 28166 17048 28172 17060
rect 28127 17020 28172 17048
rect 28166 17008 28172 17020
rect 28224 17008 28230 17060
rect 1104 16890 28888 16912
rect 1104 16838 10243 16890
rect 10295 16838 10307 16890
rect 10359 16838 10371 16890
rect 10423 16838 10435 16890
rect 10487 16838 19504 16890
rect 19556 16838 19568 16890
rect 19620 16838 19632 16890
rect 19684 16838 19696 16890
rect 19748 16838 28888 16890
rect 1104 16816 28888 16838
rect 1104 16346 28888 16368
rect 1104 16294 5612 16346
rect 5664 16294 5676 16346
rect 5728 16294 5740 16346
rect 5792 16294 5804 16346
rect 5856 16294 14874 16346
rect 14926 16294 14938 16346
rect 14990 16294 15002 16346
rect 15054 16294 15066 16346
rect 15118 16294 24135 16346
rect 24187 16294 24199 16346
rect 24251 16294 24263 16346
rect 24315 16294 24327 16346
rect 24379 16294 28888 16346
rect 1104 16272 28888 16294
rect 1104 15802 28888 15824
rect 1104 15750 10243 15802
rect 10295 15750 10307 15802
rect 10359 15750 10371 15802
rect 10423 15750 10435 15802
rect 10487 15750 19504 15802
rect 19556 15750 19568 15802
rect 19620 15750 19632 15802
rect 19684 15750 19696 15802
rect 19748 15750 28888 15802
rect 1104 15728 28888 15750
rect 14734 15512 14740 15564
rect 14792 15552 14798 15564
rect 14921 15555 14979 15561
rect 14921 15552 14933 15555
rect 14792 15524 14933 15552
rect 14792 15512 14798 15524
rect 14921 15521 14933 15524
rect 14967 15521 14979 15555
rect 14921 15515 14979 15521
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14829 15351 14887 15357
rect 14829 15348 14841 15351
rect 13872 15320 14841 15348
rect 13872 15308 13878 15320
rect 14829 15317 14841 15320
rect 14875 15317 14887 15351
rect 14829 15311 14887 15317
rect 1104 15258 28888 15280
rect 1104 15206 5612 15258
rect 5664 15206 5676 15258
rect 5728 15206 5740 15258
rect 5792 15206 5804 15258
rect 5856 15206 14874 15258
rect 14926 15206 14938 15258
rect 14990 15206 15002 15258
rect 15054 15206 15066 15258
rect 15118 15206 24135 15258
rect 24187 15206 24199 15258
rect 24251 15206 24263 15258
rect 24315 15206 24327 15258
rect 24379 15206 28888 15258
rect 1104 15184 28888 15206
rect 1578 14968 1584 15020
rect 1636 15008 1642 15020
rect 1636 14980 13124 15008
rect 1636 14968 1642 14980
rect 1394 14940 1400 14952
rect 1355 14912 1400 14940
rect 1394 14900 1400 14912
rect 1452 14900 1458 14952
rect 12250 14900 12256 14952
rect 12308 14940 12314 14952
rect 12345 14943 12403 14949
rect 12345 14940 12357 14943
rect 12308 14912 12357 14940
rect 12308 14900 12314 14912
rect 12345 14909 12357 14912
rect 12391 14909 12403 14943
rect 12345 14903 12403 14909
rect 12805 14943 12863 14949
rect 12805 14909 12817 14943
rect 12851 14940 12863 14943
rect 12894 14940 12900 14952
rect 12851 14912 12900 14940
rect 12851 14909 12863 14912
rect 12805 14903 12863 14909
rect 12820 14872 12848 14903
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 13096 14949 13124 14980
rect 12989 14943 13047 14949
rect 12989 14909 13001 14943
rect 13035 14909 13047 14943
rect 12989 14903 13047 14909
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14909 13139 14943
rect 13081 14903 13139 14909
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 13814 14940 13820 14952
rect 13219 14912 13820 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 12268 14844 12848 14872
rect 1581 14807 1639 14813
rect 1581 14773 1593 14807
rect 1627 14804 1639 14807
rect 8478 14804 8484 14816
rect 1627 14776 8484 14804
rect 1627 14773 1639 14776
rect 1581 14767 1639 14773
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 12268 14813 12296 14844
rect 12253 14807 12311 14813
rect 12253 14773 12265 14807
rect 12299 14773 12311 14807
rect 12253 14767 12311 14773
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 13004 14804 13032 14903
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 12860 14776 13032 14804
rect 13449 14807 13507 14813
rect 12860 14764 12866 14776
rect 13449 14773 13461 14807
rect 13495 14804 13507 14807
rect 13722 14804 13728 14816
rect 13495 14776 13728 14804
rect 13495 14773 13507 14776
rect 13449 14767 13507 14773
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 1104 14714 28888 14736
rect 1104 14662 10243 14714
rect 10295 14662 10307 14714
rect 10359 14662 10371 14714
rect 10423 14662 10435 14714
rect 10487 14662 19504 14714
rect 19556 14662 19568 14714
rect 19620 14662 19632 14714
rect 19684 14662 19696 14714
rect 19748 14662 28888 14714
rect 1104 14640 28888 14662
rect 8478 14492 8484 14544
rect 8536 14532 8542 14544
rect 8536 14504 12940 14532
rect 8536 14492 8542 14504
rect 12161 14467 12219 14473
rect 12161 14464 12173 14467
rect 11900 14436 12173 14464
rect 11900 14328 11928 14436
rect 12161 14433 12173 14436
rect 12207 14433 12219 14467
rect 12161 14427 12219 14433
rect 12250 14424 12256 14476
rect 12308 14464 12314 14476
rect 12621 14467 12679 14473
rect 12621 14464 12633 14467
rect 12308 14436 12633 14464
rect 12308 14424 12314 14436
rect 12621 14433 12633 14436
rect 12667 14433 12679 14467
rect 12802 14464 12808 14476
rect 12763 14436 12808 14464
rect 12621 14427 12679 14433
rect 12802 14424 12808 14436
rect 12860 14424 12866 14476
rect 12912 14473 12940 14504
rect 12897 14467 12955 14473
rect 12897 14433 12909 14467
rect 12943 14433 12955 14467
rect 12897 14427 12955 14433
rect 12989 14467 13047 14473
rect 12989 14433 13001 14467
rect 13035 14464 13047 14467
rect 13814 14464 13820 14476
rect 13035 14436 13820 14464
rect 13035 14433 13047 14436
rect 12989 14427 13047 14433
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 12066 14396 12072 14408
rect 11979 14368 12072 14396
rect 12066 14356 12072 14368
rect 12124 14396 12130 14408
rect 12820 14396 12848 14424
rect 12124 14368 12848 14396
rect 12124 14356 12130 14368
rect 13078 14328 13084 14340
rect 11900 14300 13084 14328
rect 13078 14288 13084 14300
rect 13136 14288 13142 14340
rect 13265 14263 13323 14269
rect 13265 14229 13277 14263
rect 13311 14260 13323 14263
rect 13538 14260 13544 14272
rect 13311 14232 13544 14260
rect 13311 14229 13323 14232
rect 13265 14223 13323 14229
rect 13538 14220 13544 14232
rect 13596 14220 13602 14272
rect 1104 14170 28888 14192
rect 1104 14118 5612 14170
rect 5664 14118 5676 14170
rect 5728 14118 5740 14170
rect 5792 14118 5804 14170
rect 5856 14118 14874 14170
rect 14926 14118 14938 14170
rect 14990 14118 15002 14170
rect 15054 14118 15066 14170
rect 15118 14118 24135 14170
rect 24187 14118 24199 14170
rect 24251 14118 24263 14170
rect 24315 14118 24327 14170
rect 24379 14118 28888 14170
rect 1104 14096 28888 14118
rect 12066 13988 12072 14000
rect 10980 13960 12072 13988
rect 10980 13861 11008 13960
rect 12066 13948 12072 13960
rect 12124 13948 12130 14000
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13920 11115 13923
rect 11103 13892 12480 13920
rect 11103 13889 11115 13892
rect 11057 13883 11115 13889
rect 10965 13855 11023 13861
rect 10965 13821 10977 13855
rect 11011 13821 11023 13855
rect 10965 13815 11023 13821
rect 11149 13855 11207 13861
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 12452 13852 12480 13892
rect 13170 13852 13176 13864
rect 13228 13861 13234 13864
rect 11195 13824 12388 13852
rect 12452 13824 13176 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 12360 13784 12388 13824
rect 13170 13812 13176 13824
rect 13228 13815 13240 13861
rect 13446 13852 13452 13864
rect 13407 13824 13452 13852
rect 13228 13812 13234 13815
rect 13446 13812 13452 13824
rect 13504 13852 13510 13864
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13504 13824 13921 13852
rect 13504 13812 13510 13824
rect 13909 13821 13921 13824
rect 13955 13821 13967 13855
rect 27982 13852 27988 13864
rect 13909 13815 13967 13821
rect 16546 13824 27988 13852
rect 12894 13784 12900 13796
rect 12360 13756 12900 13784
rect 12894 13744 12900 13756
rect 12952 13744 12958 13796
rect 14176 13787 14234 13793
rect 14176 13753 14188 13787
rect 14222 13784 14234 13787
rect 14366 13784 14372 13796
rect 14222 13756 14372 13784
rect 14222 13753 14234 13756
rect 14176 13747 14234 13753
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 12069 13719 12127 13725
rect 12069 13685 12081 13719
rect 12115 13716 12127 13719
rect 12158 13716 12164 13728
rect 12115 13688 12164 13716
rect 12115 13685 12127 13688
rect 12069 13679 12127 13685
rect 12158 13676 12164 13688
rect 12216 13676 12222 13728
rect 15286 13716 15292 13728
rect 15247 13688 15292 13716
rect 15286 13676 15292 13688
rect 15344 13716 15350 13728
rect 16546 13716 16574 13824
rect 27982 13812 27988 13824
rect 28040 13812 28046 13864
rect 15344 13688 16574 13716
rect 15344 13676 15350 13688
rect 1104 13626 28888 13648
rect 1104 13574 10243 13626
rect 10295 13574 10307 13626
rect 10359 13574 10371 13626
rect 10423 13574 10435 13626
rect 10487 13574 19504 13626
rect 19556 13574 19568 13626
rect 19620 13574 19632 13626
rect 19684 13574 19696 13626
rect 19748 13574 28888 13626
rect 1104 13552 28888 13574
rect 11701 13515 11759 13521
rect 11701 13481 11713 13515
rect 11747 13512 11759 13515
rect 12250 13512 12256 13524
rect 11747 13484 12256 13512
rect 11747 13481 11759 13484
rect 11701 13475 11759 13481
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 1578 13336 1584 13388
rect 1636 13376 1642 13388
rect 10781 13379 10839 13385
rect 10781 13376 10793 13379
rect 1636 13348 10793 13376
rect 1636 13336 1642 13348
rect 10781 13345 10793 13348
rect 10827 13345 10839 13379
rect 10781 13339 10839 13345
rect 10873 13379 10931 13385
rect 10873 13345 10885 13379
rect 10919 13376 10931 13379
rect 11977 13379 12035 13385
rect 11977 13376 11989 13379
rect 10919 13348 11989 13376
rect 10919 13345 10931 13348
rect 10873 13339 10931 13345
rect 11977 13345 11989 13348
rect 12023 13345 12035 13379
rect 12158 13376 12164 13388
rect 12119 13348 12164 13376
rect 11977 13339 12035 13345
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 12894 13336 12900 13388
rect 12952 13376 12958 13388
rect 13265 13379 13323 13385
rect 13265 13376 13277 13379
rect 12952 13348 13277 13376
rect 12952 13336 12958 13348
rect 13265 13345 13277 13348
rect 13311 13345 13323 13379
rect 13265 13339 13323 13345
rect 13449 13379 13507 13385
rect 13449 13345 13461 13379
rect 13495 13376 13507 13379
rect 15286 13376 15292 13388
rect 13495 13348 15292 13376
rect 13495 13345 13507 13348
rect 13449 13339 13507 13345
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 9824 13280 11897 13308
rect 9824 13268 9830 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 12066 13308 12072 13320
rect 12027 13280 12072 13308
rect 11885 13271 11943 13277
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 13136 13280 13185 13308
rect 13136 13268 13142 13280
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13633 13175 13691 13181
rect 13633 13141 13645 13175
rect 13679 13172 13691 13175
rect 13998 13172 14004 13184
rect 13679 13144 14004 13172
rect 13679 13141 13691 13144
rect 13633 13135 13691 13141
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 1104 13082 28888 13104
rect 1104 13030 5612 13082
rect 5664 13030 5676 13082
rect 5728 13030 5740 13082
rect 5792 13030 5804 13082
rect 5856 13030 14874 13082
rect 14926 13030 14938 13082
rect 14990 13030 15002 13082
rect 15054 13030 15066 13082
rect 15118 13030 24135 13082
rect 24187 13030 24199 13082
rect 24251 13030 24263 13082
rect 24315 13030 24327 13082
rect 24379 13030 28888 13082
rect 1104 13008 28888 13030
rect 13078 12928 13084 12980
rect 13136 12968 13142 12980
rect 13541 12971 13599 12977
rect 13541 12968 13553 12971
rect 13136 12940 13553 12968
rect 13136 12928 13142 12940
rect 13541 12937 13553 12940
rect 13587 12937 13599 12971
rect 14366 12968 14372 12980
rect 14327 12940 14372 12968
rect 13541 12931 13599 12937
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 10962 12764 10968 12776
rect 10008 12736 10968 12764
rect 10008 12724 10014 12736
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 12158 12764 12164 12776
rect 12119 12736 12164 12764
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 13998 12764 14004 12776
rect 13959 12736 14004 12764
rect 13998 12724 14004 12736
rect 14056 12724 14062 12776
rect 12428 12699 12486 12705
rect 12428 12665 12440 12699
rect 12474 12696 12486 12699
rect 12618 12696 12624 12708
rect 12474 12668 12624 12696
rect 12474 12665 12486 12668
rect 12428 12659 12486 12665
rect 12618 12656 12624 12668
rect 12676 12656 12682 12708
rect 14185 12699 14243 12705
rect 14185 12665 14197 12699
rect 14231 12696 14243 12699
rect 14550 12696 14556 12708
rect 14231 12668 14556 12696
rect 14231 12665 14243 12668
rect 14185 12659 14243 12665
rect 14550 12656 14556 12668
rect 14608 12656 14614 12708
rect 11057 12631 11115 12637
rect 11057 12597 11069 12631
rect 11103 12628 11115 12631
rect 12526 12628 12532 12640
rect 11103 12600 12532 12628
rect 11103 12597 11115 12600
rect 11057 12591 11115 12597
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 1104 12538 28888 12560
rect 1104 12486 10243 12538
rect 10295 12486 10307 12538
rect 10359 12486 10371 12538
rect 10423 12486 10435 12538
rect 10487 12486 19504 12538
rect 19556 12486 19568 12538
rect 19620 12486 19632 12538
rect 19684 12486 19696 12538
rect 19748 12486 28888 12538
rect 1104 12464 28888 12486
rect 12618 12424 12624 12436
rect 12579 12396 12624 12424
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 13354 12384 13360 12436
rect 13412 12424 13418 12436
rect 13722 12424 13728 12436
rect 13412 12396 13728 12424
rect 13412 12384 13418 12396
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 12158 12356 12164 12368
rect 10244 12328 12164 12356
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 10244 12229 10272 12328
rect 12158 12316 12164 12328
rect 12216 12356 12222 12368
rect 13446 12356 13452 12368
rect 12216 12328 13452 12356
rect 12216 12316 12222 12328
rect 13446 12316 13452 12328
rect 13504 12316 13510 12368
rect 14458 12316 14464 12368
rect 14516 12356 14522 12368
rect 14516 12328 14964 12356
rect 14516 12316 14522 12328
rect 10496 12291 10554 12297
rect 10496 12257 10508 12291
rect 10542 12288 10554 12291
rect 11514 12288 11520 12300
rect 10542 12260 11520 12288
rect 10542 12257 10554 12260
rect 10496 12251 10554 12257
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 12805 12291 12863 12297
rect 12805 12288 12817 12291
rect 12728 12260 12817 12288
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 9824 12192 10241 12220
rect 9824 12180 9830 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 12728 12152 12756 12260
rect 12805 12257 12817 12260
rect 12851 12257 12863 12291
rect 12805 12251 12863 12257
rect 13081 12291 13139 12297
rect 13081 12257 13093 12291
rect 13127 12288 13139 12291
rect 13170 12288 13176 12300
rect 13127 12260 13176 12288
rect 13127 12257 13139 12260
rect 13081 12251 13139 12257
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 13722 12288 13728 12300
rect 13679 12260 13728 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 14936 12297 14964 12328
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12257 14795 12291
rect 14737 12251 14795 12257
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 12894 12220 12900 12232
rect 12855 12192 12900 12220
rect 12894 12180 12900 12192
rect 12952 12180 12958 12232
rect 12986 12180 12992 12232
rect 13044 12220 13050 12232
rect 14752 12220 14780 12251
rect 15562 12220 15568 12232
rect 13044 12192 13089 12220
rect 14752 12192 15568 12220
rect 13044 12180 13050 12192
rect 15562 12180 15568 12192
rect 15620 12180 15626 12232
rect 13262 12152 13268 12164
rect 12728 12124 13268 12152
rect 13262 12112 13268 12124
rect 13320 12112 13326 12164
rect 11609 12087 11667 12093
rect 11609 12053 11621 12087
rect 11655 12084 11667 12087
rect 12434 12084 12440 12096
rect 11655 12056 12440 12084
rect 11655 12053 11667 12056
rect 11609 12047 11667 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 13817 12087 13875 12093
rect 13817 12084 13829 12087
rect 13504 12056 13829 12084
rect 13504 12044 13510 12056
rect 13817 12053 13829 12056
rect 13863 12084 13875 12087
rect 14550 12084 14556 12096
rect 13863 12056 14556 12084
rect 13863 12053 13875 12056
rect 13817 12047 13875 12053
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 14642 12044 14648 12096
rect 14700 12084 14706 12096
rect 14921 12087 14979 12093
rect 14921 12084 14933 12087
rect 14700 12056 14933 12084
rect 14700 12044 14706 12056
rect 14921 12053 14933 12056
rect 14967 12053 14979 12087
rect 14921 12047 14979 12053
rect 1104 11994 28888 12016
rect 1104 11942 5612 11994
rect 5664 11942 5676 11994
rect 5728 11942 5740 11994
rect 5792 11942 5804 11994
rect 5856 11942 14874 11994
rect 14926 11942 14938 11994
rect 14990 11942 15002 11994
rect 15054 11942 15066 11994
rect 15118 11942 24135 11994
rect 24187 11942 24199 11994
rect 24251 11942 24263 11994
rect 24315 11942 24327 11994
rect 24379 11942 28888 11994
rect 1104 11920 28888 11942
rect 12805 11883 12863 11889
rect 12805 11849 12817 11883
rect 12851 11880 12863 11883
rect 12894 11880 12900 11892
rect 12851 11852 12900 11880
rect 12851 11849 12863 11852
rect 12805 11843 12863 11849
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 13262 11880 13268 11892
rect 13223 11852 13268 11880
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 13633 11883 13691 11889
rect 13633 11849 13645 11883
rect 13679 11880 13691 11883
rect 14090 11880 14096 11892
rect 13679 11852 14096 11880
rect 13679 11849 13691 11852
rect 13633 11843 13691 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 9769 11815 9827 11821
rect 9769 11781 9781 11815
rect 9815 11812 9827 11815
rect 11054 11812 11060 11824
rect 9815 11784 11060 11812
rect 9815 11781 9827 11784
rect 9769 11775 9827 11781
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 12345 11747 12403 11753
rect 12345 11744 12357 11747
rect 9876 11716 12357 11744
rect 9876 11685 9904 11716
rect 12345 11713 12357 11716
rect 12391 11744 12403 11747
rect 12710 11744 12716 11756
rect 12391 11716 12716 11744
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11744 14979 11747
rect 15102 11744 15108 11756
rect 14967 11716 15108 11744
rect 14967 11713 14979 11716
rect 14921 11707 14979 11713
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 9861 11679 9919 11685
rect 9861 11645 9873 11679
rect 9907 11645 9919 11679
rect 9861 11639 9919 11645
rect 10321 11679 10379 11685
rect 10321 11645 10333 11679
rect 10367 11645 10379 11679
rect 10321 11639 10379 11645
rect 10505 11679 10563 11685
rect 10505 11645 10517 11679
rect 10551 11676 10563 11679
rect 10870 11676 10876 11688
rect 10551 11648 10876 11676
rect 10551 11645 10563 11648
rect 10505 11639 10563 11645
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 10336 11608 10364 11639
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 10962 11636 10968 11688
rect 11020 11676 11026 11688
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11020 11648 12081 11676
rect 11020 11636 11026 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12250 11676 12256 11688
rect 12211 11648 12256 11676
rect 12069 11639 12127 11645
rect 12250 11636 12256 11648
rect 12308 11636 12314 11688
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 12621 11679 12679 11685
rect 12621 11645 12633 11679
rect 12667 11676 12679 11679
rect 13078 11676 13084 11688
rect 12667 11648 13084 11676
rect 12667 11645 12679 11648
rect 12621 11639 12679 11645
rect 9732 11580 10364 11608
rect 12452 11608 12480 11639
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 13354 11636 13360 11688
rect 13412 11676 13418 11688
rect 13449 11679 13507 11685
rect 13449 11676 13461 11679
rect 13412 11648 13461 11676
rect 13412 11636 13418 11648
rect 13449 11645 13461 11648
rect 13495 11645 13507 11679
rect 13630 11676 13636 11688
rect 13591 11648 13636 11676
rect 13449 11639 13507 11645
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 14642 11676 14648 11688
rect 14603 11648 14648 11676
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 15657 11679 15715 11685
rect 15657 11645 15669 11679
rect 15703 11676 15715 11679
rect 16114 11676 16120 11688
rect 15703 11648 16120 11676
rect 15703 11645 15715 11648
rect 15657 11639 15715 11645
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 14458 11608 14464 11620
rect 12452 11580 14464 11608
rect 9732 11568 9738 11580
rect 14458 11568 14464 11580
rect 14516 11568 14522 11620
rect 10686 11540 10692 11552
rect 10647 11512 10692 11540
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 14274 11540 14280 11552
rect 14235 11512 14280 11540
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 14737 11543 14795 11549
rect 14737 11509 14749 11543
rect 14783 11540 14795 11543
rect 15562 11540 15568 11552
rect 14783 11512 15568 11540
rect 14783 11509 14795 11512
rect 14737 11503 14795 11509
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 1104 11450 28888 11472
rect 1104 11398 10243 11450
rect 10295 11398 10307 11450
rect 10359 11398 10371 11450
rect 10423 11398 10435 11450
rect 10487 11398 19504 11450
rect 19556 11398 19568 11450
rect 19620 11398 19632 11450
rect 19684 11398 19696 11450
rect 19748 11398 28888 11450
rect 1104 11376 28888 11398
rect 11514 11336 11520 11348
rect 11475 11308 11520 11336
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 12710 11336 12716 11348
rect 12671 11308 12716 11336
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13541 11339 13599 11345
rect 13541 11336 13553 11339
rect 13044 11308 13553 11336
rect 13044 11296 13050 11308
rect 13541 11305 13553 11308
rect 13587 11305 13599 11339
rect 16114 11336 16120 11348
rect 16075 11308 16120 11336
rect 13541 11299 13599 11305
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 10790 11271 10848 11277
rect 10790 11268 10802 11271
rect 10744 11240 10802 11268
rect 10744 11228 10750 11240
rect 10790 11237 10802 11240
rect 10836 11237 10848 11271
rect 10790 11231 10848 11237
rect 10962 11228 10968 11280
rect 11020 11268 11026 11280
rect 12434 11268 12440 11280
rect 11020 11240 11744 11268
rect 11020 11228 11026 11240
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 11716 11209 11744 11240
rect 11900 11240 12440 11268
rect 11900 11209 11928 11240
rect 12434 11228 12440 11240
rect 12492 11268 12498 11280
rect 12529 11271 12587 11277
rect 12529 11268 12541 11271
rect 12492 11240 12541 11268
rect 12492 11228 12498 11240
rect 12529 11237 12541 11240
rect 12575 11237 12587 11271
rect 12529 11231 12587 11237
rect 14642 11228 14648 11280
rect 14700 11268 14706 11280
rect 14982 11271 15040 11277
rect 14982 11268 14994 11271
rect 14700 11240 14994 11268
rect 14700 11228 14706 11240
rect 14982 11237 14994 11240
rect 15028 11237 15040 11271
rect 14982 11231 15040 11237
rect 11057 11203 11115 11209
rect 11057 11200 11069 11203
rect 9824 11172 11069 11200
rect 9824 11160 9830 11172
rect 11057 11169 11069 11172
rect 11103 11169 11115 11203
rect 11057 11163 11115 11169
rect 11701 11203 11759 11209
rect 11701 11169 11713 11203
rect 11747 11169 11759 11203
rect 11701 11163 11759 11169
rect 11885 11203 11943 11209
rect 11885 11169 11897 11203
rect 11931 11169 11943 11203
rect 11885 11163 11943 11169
rect 11716 11132 11744 11163
rect 11974 11160 11980 11212
rect 12032 11200 12038 11212
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 12032 11172 12357 11200
rect 12032 11160 12038 11172
rect 12345 11169 12357 11172
rect 12391 11169 12403 11203
rect 12345 11163 12403 11169
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11169 13691 11203
rect 13814 11200 13820 11212
rect 13775 11172 13820 11200
rect 13633 11163 13691 11169
rect 13538 11132 13544 11144
rect 11716 11104 13544 11132
rect 12360 11076 12388 11104
rect 13538 11092 13544 11104
rect 13596 11092 13602 11144
rect 13648 11132 13676 11163
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 14550 11160 14556 11212
rect 14608 11200 14614 11212
rect 14737 11203 14795 11209
rect 14737 11200 14749 11203
rect 14608 11172 14749 11200
rect 14608 11160 14614 11172
rect 14737 11169 14749 11172
rect 14783 11169 14795 11203
rect 14737 11163 14795 11169
rect 14642 11132 14648 11144
rect 13648 11104 14648 11132
rect 14642 11092 14648 11104
rect 14700 11092 14706 11144
rect 12342 11024 12348 11076
rect 12400 11024 12406 11076
rect 9674 10996 9680 11008
rect 9635 10968 9680 10996
rect 9674 10956 9680 10968
rect 9732 10956 9738 11008
rect 13354 10996 13360 11008
rect 13315 10968 13360 10996
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 1104 10906 28888 10928
rect 1104 10854 5612 10906
rect 5664 10854 5676 10906
rect 5728 10854 5740 10906
rect 5792 10854 5804 10906
rect 5856 10854 14874 10906
rect 14926 10854 14938 10906
rect 14990 10854 15002 10906
rect 15054 10854 15066 10906
rect 15118 10854 24135 10906
rect 24187 10854 24199 10906
rect 24251 10854 24263 10906
rect 24315 10854 24327 10906
rect 24379 10854 28888 10906
rect 1104 10832 28888 10854
rect 9950 10792 9956 10804
rect 9911 10764 9956 10792
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 10962 10792 10968 10804
rect 10923 10764 10968 10792
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 11149 10795 11207 10801
rect 11149 10761 11161 10795
rect 11195 10792 11207 10795
rect 12250 10792 12256 10804
rect 11195 10764 12256 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 12250 10752 12256 10764
rect 12308 10792 12314 10804
rect 12345 10795 12403 10801
rect 12345 10792 12357 10795
rect 12308 10764 12357 10792
rect 12308 10752 12314 10764
rect 12345 10761 12357 10764
rect 12391 10761 12403 10795
rect 12526 10792 12532 10804
rect 12487 10764 12532 10792
rect 12345 10755 12403 10761
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 12805 10795 12863 10801
rect 12805 10761 12817 10795
rect 12851 10792 12863 10795
rect 13354 10792 13360 10804
rect 12851 10764 13360 10792
rect 12851 10761 12863 10764
rect 12805 10755 12863 10761
rect 13354 10752 13360 10764
rect 13412 10752 13418 10804
rect 13449 10795 13507 10801
rect 13449 10761 13461 10795
rect 13495 10792 13507 10795
rect 13814 10792 13820 10804
rect 13495 10764 13820 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 13814 10752 13820 10764
rect 13872 10752 13878 10804
rect 14274 10792 14280 10804
rect 14235 10764 14280 10792
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 14642 10752 14648 10804
rect 14700 10792 14706 10804
rect 15749 10795 15807 10801
rect 15749 10792 15761 10795
rect 14700 10764 15761 10792
rect 14700 10752 14706 10764
rect 15749 10761 15761 10764
rect 15795 10761 15807 10795
rect 15749 10755 15807 10761
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10761 15991 10795
rect 15933 10755 15991 10761
rect 11054 10684 11060 10736
rect 11112 10724 11118 10736
rect 12437 10727 12495 10733
rect 12437 10724 12449 10727
rect 11112 10696 12449 10724
rect 11112 10684 11118 10696
rect 12437 10693 12449 10696
rect 12483 10693 12495 10727
rect 12437 10687 12495 10693
rect 13280 10696 15332 10724
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 10137 10591 10195 10597
rect 10137 10588 10149 10591
rect 9732 10560 10149 10588
rect 9732 10548 9738 10560
rect 10137 10557 10149 10560
rect 10183 10588 10195 10591
rect 10183 10560 10824 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 10321 10523 10379 10529
rect 10321 10489 10333 10523
rect 10367 10520 10379 10523
rect 10594 10520 10600 10532
rect 10367 10492 10600 10520
rect 10367 10489 10379 10492
rect 10321 10483 10379 10489
rect 10594 10480 10600 10492
rect 10652 10480 10658 10532
rect 10796 10529 10824 10560
rect 11514 10548 11520 10600
rect 11572 10588 11578 10600
rect 13280 10597 13308 10696
rect 13538 10616 13544 10668
rect 13596 10656 13602 10668
rect 15304 10665 15332 10696
rect 15378 10684 15384 10736
rect 15436 10724 15442 10736
rect 15948 10724 15976 10755
rect 15436 10696 15976 10724
rect 15436 10684 15442 10696
rect 15289 10659 15347 10665
rect 13596 10628 15148 10656
rect 13596 10616 13602 10628
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 11572 10560 12081 10588
rect 11572 10548 11578 10560
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 13265 10591 13323 10597
rect 13265 10557 13277 10591
rect 13311 10557 13323 10591
rect 13265 10551 13323 10557
rect 13449 10591 13507 10597
rect 13449 10557 13461 10591
rect 13495 10557 13507 10591
rect 13449 10551 13507 10557
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10588 13967 10591
rect 14182 10588 14188 10600
rect 13955 10560 14188 10588
rect 13955 10557 13967 10560
rect 13909 10551 13967 10557
rect 10781 10523 10839 10529
rect 10781 10489 10793 10523
rect 10827 10489 10839 10523
rect 10781 10483 10839 10489
rect 10962 10412 10968 10464
rect 11020 10461 11026 10464
rect 11020 10455 11044 10461
rect 11032 10421 11044 10455
rect 12158 10452 12164 10464
rect 12119 10424 12164 10452
rect 11020 10415 11044 10421
rect 11020 10412 11026 10415
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 13464 10452 13492 10551
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 15120 10597 15148 10628
rect 15289 10625 15301 10659
rect 15335 10656 15347 10659
rect 16114 10656 16120 10668
rect 15335 10628 16120 10656
rect 15335 10625 15347 10628
rect 15289 10619 15347 10625
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 14277 10591 14335 10597
rect 14277 10557 14289 10591
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 15105 10591 15163 10597
rect 15105 10557 15117 10591
rect 15151 10557 15163 10591
rect 15105 10551 15163 10557
rect 13814 10480 13820 10532
rect 13872 10520 13878 10532
rect 14292 10520 14320 10551
rect 13872 10492 14320 10520
rect 13872 10480 13878 10492
rect 14366 10480 14372 10532
rect 14424 10520 14430 10532
rect 14424 10492 15056 10520
rect 14424 10480 14430 10492
rect 13906 10452 13912 10464
rect 13464 10424 13912 10452
rect 13906 10412 13912 10424
rect 13964 10412 13970 10464
rect 14090 10452 14096 10464
rect 14051 10424 14096 10452
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 14240 10424 14933 10452
rect 14240 10412 14246 10424
rect 14921 10421 14933 10424
rect 14967 10421 14979 10455
rect 15028 10452 15056 10492
rect 15562 10480 15568 10532
rect 15620 10520 15626 10532
rect 16117 10523 16175 10529
rect 16117 10520 16129 10523
rect 15620 10492 16129 10520
rect 15620 10480 15626 10492
rect 16117 10489 16129 10492
rect 16163 10489 16175 10523
rect 16117 10483 16175 10489
rect 15912 10455 15970 10461
rect 15912 10452 15924 10455
rect 15028 10424 15924 10452
rect 14921 10415 14979 10421
rect 15912 10421 15924 10424
rect 15958 10421 15970 10455
rect 15912 10415 15970 10421
rect 1104 10362 28888 10384
rect 1104 10310 10243 10362
rect 10295 10310 10307 10362
rect 10359 10310 10371 10362
rect 10423 10310 10435 10362
rect 10487 10310 19504 10362
rect 19556 10310 19568 10362
rect 19620 10310 19632 10362
rect 19684 10310 19696 10362
rect 19748 10310 28888 10362
rect 1104 10288 28888 10310
rect 10594 10208 10600 10260
rect 10652 10248 10658 10260
rect 13081 10251 13139 10257
rect 13081 10248 13093 10251
rect 10652 10220 13093 10248
rect 10652 10208 10658 10220
rect 13081 10217 13093 10220
rect 13127 10217 13139 10251
rect 16114 10248 16120 10260
rect 16075 10220 16120 10248
rect 13081 10211 13139 10217
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 10962 10140 10968 10192
rect 11020 10180 11026 10192
rect 12713 10183 12771 10189
rect 12713 10180 12725 10183
rect 11020 10152 12725 10180
rect 11020 10140 11026 10152
rect 12713 10149 12725 10152
rect 12759 10149 12771 10183
rect 12713 10143 12771 10149
rect 10134 10072 10140 10124
rect 10192 10112 10198 10124
rect 10301 10115 10359 10121
rect 10301 10112 10313 10115
rect 10192 10084 10313 10112
rect 10192 10072 10198 10084
rect 10301 10081 10313 10084
rect 10347 10081 10359 10115
rect 10301 10075 10359 10081
rect 11974 10072 11980 10124
rect 12032 10112 12038 10124
rect 12069 10115 12127 10121
rect 12069 10112 12081 10115
rect 12032 10084 12081 10112
rect 12032 10072 12038 10084
rect 12069 10081 12081 10084
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 10045 10047 10103 10053
rect 10045 10044 10057 10047
rect 9824 10016 10057 10044
rect 9824 10004 9830 10016
rect 10045 10013 10057 10016
rect 10091 10013 10103 10047
rect 12084 10044 12112 10075
rect 12158 10072 12164 10124
rect 12216 10112 12222 10124
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 12216 10084 12265 10112
rect 12216 10072 12222 10084
rect 12253 10081 12265 10084
rect 12299 10081 12311 10115
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 12253 10075 12311 10081
rect 12406 10084 12909 10112
rect 12406 10044 12434 10084
rect 12897 10081 12909 10084
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 13633 10115 13691 10121
rect 13633 10081 13645 10115
rect 13679 10112 13691 10115
rect 14182 10112 14188 10124
rect 13679 10084 14188 10112
rect 13679 10081 13691 10084
rect 13633 10075 13691 10081
rect 14182 10072 14188 10084
rect 14240 10072 14246 10124
rect 14993 10115 15051 10121
rect 14993 10112 15005 10115
rect 14292 10084 15005 10112
rect 12084 10016 12434 10044
rect 10045 10007 10103 10013
rect 13814 9976 13820 9988
rect 13727 9948 13820 9976
rect 13814 9936 13820 9948
rect 13872 9976 13878 9988
rect 14292 9976 14320 10084
rect 14993 10081 15005 10084
rect 15039 10081 15051 10115
rect 14993 10075 15051 10081
rect 14642 10004 14648 10056
rect 14700 10044 14706 10056
rect 14737 10047 14795 10053
rect 14737 10044 14749 10047
rect 14700 10016 14749 10044
rect 14700 10004 14706 10016
rect 14737 10013 14749 10016
rect 14783 10013 14795 10047
rect 14737 10007 14795 10013
rect 13872 9948 14320 9976
rect 13872 9936 13878 9948
rect 11422 9908 11428 9920
rect 11383 9880 11428 9908
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 11882 9908 11888 9920
rect 11843 9880 11888 9908
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 1104 9818 28888 9840
rect 1104 9766 5612 9818
rect 5664 9766 5676 9818
rect 5728 9766 5740 9818
rect 5792 9766 5804 9818
rect 5856 9766 14874 9818
rect 14926 9766 14938 9818
rect 14990 9766 15002 9818
rect 15054 9766 15066 9818
rect 15118 9766 24135 9818
rect 24187 9766 24199 9818
rect 24251 9766 24263 9818
rect 24315 9766 24327 9818
rect 24379 9766 28888 9818
rect 1104 9744 28888 9766
rect 12158 9704 12164 9716
rect 12119 9676 12164 9704
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 13909 9707 13967 9713
rect 13909 9673 13921 9707
rect 13955 9704 13967 9707
rect 14274 9704 14280 9716
rect 13955 9676 14280 9704
rect 13955 9673 13967 9676
rect 13909 9667 13967 9673
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 14476 9608 16068 9636
rect 9766 9568 9772 9580
rect 9727 9540 9772 9568
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 12069 9571 12127 9577
rect 12069 9568 12081 9571
rect 11572 9540 12081 9568
rect 11572 9528 11578 9540
rect 12069 9537 12081 9540
rect 12115 9537 12127 9571
rect 12069 9531 12127 9537
rect 13906 9528 13912 9580
rect 13964 9568 13970 9580
rect 14476 9577 14504 9608
rect 14461 9571 14519 9577
rect 14461 9568 14473 9571
rect 13964 9540 14473 9568
rect 13964 9528 13970 9540
rect 14461 9537 14473 9540
rect 14507 9537 14519 9571
rect 15286 9568 15292 9580
rect 15247 9540 15292 9568
rect 14461 9531 14519 9537
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 12250 9500 12256 9512
rect 12211 9472 12256 9500
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 12345 9503 12403 9509
rect 12345 9469 12357 9503
rect 12391 9469 12403 9503
rect 13814 9500 13820 9512
rect 13775 9472 13820 9500
rect 12345 9463 12403 9469
rect 10036 9435 10094 9441
rect 10036 9401 10048 9435
rect 10082 9432 10094 9435
rect 10870 9432 10876 9444
rect 10082 9404 10876 9432
rect 10082 9401 10094 9404
rect 10036 9395 10094 9401
rect 10870 9392 10876 9404
rect 10928 9392 10934 9444
rect 12066 9432 12072 9444
rect 11164 9404 12072 9432
rect 11164 9373 11192 9404
rect 12066 9392 12072 9404
rect 12124 9432 12130 9444
rect 12360 9432 12388 9463
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 14001 9503 14059 9509
rect 14001 9469 14013 9503
rect 14047 9500 14059 9503
rect 14047 9472 14872 9500
rect 14047 9469 14059 9472
rect 14001 9463 14059 9469
rect 12124 9404 12388 9432
rect 12124 9392 12130 9404
rect 14458 9392 14464 9444
rect 14516 9432 14522 9444
rect 14844 9441 14872 9472
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 16040 9509 16068 9608
rect 15473 9503 15531 9509
rect 15473 9500 15485 9503
rect 15252 9472 15485 9500
rect 15252 9460 15258 9472
rect 15473 9469 15485 9472
rect 15519 9469 15531 9503
rect 15473 9463 15531 9469
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9469 15623 9503
rect 15565 9463 15623 9469
rect 16025 9503 16083 9509
rect 16025 9469 16037 9503
rect 16071 9469 16083 9503
rect 16025 9463 16083 9469
rect 14645 9435 14703 9441
rect 14645 9432 14657 9435
rect 14516 9404 14657 9432
rect 14516 9392 14522 9404
rect 14645 9401 14657 9404
rect 14691 9401 14703 9435
rect 14645 9395 14703 9401
rect 14829 9435 14887 9441
rect 14829 9401 14841 9435
rect 14875 9432 14887 9435
rect 15289 9435 15347 9441
rect 15289 9432 15301 9435
rect 14875 9404 15301 9432
rect 14875 9401 14887 9404
rect 14829 9395 14887 9401
rect 15289 9401 15301 9404
rect 15335 9401 15347 9435
rect 15580 9432 15608 9463
rect 16206 9432 16212 9444
rect 15580 9404 16212 9432
rect 15289 9395 15347 9401
rect 16206 9392 16212 9404
rect 16264 9392 16270 9444
rect 11149 9367 11207 9373
rect 11149 9333 11161 9367
rect 11195 9333 11207 9367
rect 16114 9364 16120 9376
rect 16075 9336 16120 9364
rect 11149 9327 11207 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 1104 9274 28888 9296
rect 1104 9222 10243 9274
rect 10295 9222 10307 9274
rect 10359 9222 10371 9274
rect 10423 9222 10435 9274
rect 10487 9222 19504 9274
rect 19556 9222 19568 9274
rect 19620 9222 19632 9274
rect 19684 9222 19696 9274
rect 19748 9222 28888 9274
rect 1104 9200 28888 9222
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10413 9163 10471 9169
rect 10413 9160 10425 9163
rect 10192 9132 10425 9160
rect 10192 9120 10198 9132
rect 10413 9129 10425 9132
rect 10459 9129 10471 9163
rect 10962 9160 10968 9172
rect 10923 9132 10968 9160
rect 10413 9123 10471 9129
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11149 9163 11207 9169
rect 11149 9129 11161 9163
rect 11195 9160 11207 9163
rect 11514 9160 11520 9172
rect 11195 9132 11520 9160
rect 11195 9129 11207 9132
rect 11149 9123 11207 9129
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 15004 9095 15062 9101
rect 15004 9061 15016 9095
rect 15050 9092 15062 9095
rect 16114 9092 16120 9104
rect 15050 9064 16120 9092
rect 15050 9061 15062 9064
rect 15004 9055 15062 9061
rect 16114 9052 16120 9064
rect 16172 9052 16178 9104
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 10594 9024 10600 9036
rect 10551 8996 10600 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 11146 9027 11204 9033
rect 11146 8993 11158 9027
rect 11192 9024 11204 9027
rect 11422 9024 11428 9036
rect 11192 8996 11428 9024
rect 11192 8993 11204 8996
rect 11146 8987 11204 8993
rect 11422 8984 11428 8996
rect 11480 9024 11486 9036
rect 11609 9027 11667 9033
rect 11609 9024 11621 9027
rect 11480 8996 11621 9024
rect 11480 8984 11486 8996
rect 11609 8993 11621 8996
rect 11655 8993 11667 9027
rect 11609 8987 11667 8993
rect 11790 8984 11796 9036
rect 11848 9024 11854 9036
rect 12069 9027 12127 9033
rect 12069 9024 12081 9027
rect 11848 8996 12081 9024
rect 11848 8984 11854 8996
rect 12069 8993 12081 8996
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 14642 8984 14648 9036
rect 14700 9024 14706 9036
rect 14737 9027 14795 9033
rect 14737 9024 14749 9027
rect 14700 8996 14749 9024
rect 14700 8984 14706 8996
rect 14737 8993 14749 8996
rect 14783 8993 14795 9027
rect 14737 8987 14795 8993
rect 10134 8848 10140 8900
rect 10192 8888 10198 8900
rect 13357 8891 13415 8897
rect 13357 8888 13369 8891
rect 10192 8860 13369 8888
rect 10192 8848 10198 8860
rect 13357 8857 13369 8860
rect 13403 8888 13415 8891
rect 13722 8888 13728 8900
rect 13403 8860 13728 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 13722 8848 13728 8860
rect 13780 8848 13786 8900
rect 11514 8820 11520 8832
rect 11475 8792 11520 8820
rect 11514 8780 11520 8792
rect 11572 8780 11578 8832
rect 16114 8820 16120 8832
rect 16075 8792 16120 8820
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 1104 8730 28888 8752
rect 1104 8678 5612 8730
rect 5664 8678 5676 8730
rect 5728 8678 5740 8730
rect 5792 8678 5804 8730
rect 5856 8678 14874 8730
rect 14926 8678 14938 8730
rect 14990 8678 15002 8730
rect 15054 8678 15066 8730
rect 15118 8678 24135 8730
rect 24187 8678 24199 8730
rect 24251 8678 24263 8730
rect 24315 8678 24327 8730
rect 24379 8678 28888 8730
rect 1104 8656 28888 8678
rect 10870 8616 10876 8628
rect 10831 8588 10876 8616
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 11572 8588 12173 8616
rect 11572 8576 11578 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 15286 8480 15292 8492
rect 13832 8452 15292 8480
rect 10965 8415 11023 8421
rect 10965 8381 10977 8415
rect 11011 8412 11023 8415
rect 11882 8412 11888 8424
rect 11011 8384 11888 8412
rect 11011 8381 11023 8384
rect 10965 8375 11023 8381
rect 11882 8372 11888 8384
rect 11940 8372 11946 8424
rect 12066 8412 12072 8424
rect 12027 8384 12072 8412
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 12250 8412 12256 8424
rect 12211 8384 12256 8412
rect 12250 8372 12256 8384
rect 12308 8412 12314 8424
rect 13832 8421 13860 8452
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 12308 8384 13737 8412
rect 12308 8372 12314 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 13817 8415 13875 8421
rect 13817 8381 13829 8415
rect 13863 8381 13875 8415
rect 14550 8412 14556 8424
rect 14511 8384 14556 8412
rect 13817 8375 13875 8381
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 14645 8415 14703 8421
rect 14645 8381 14657 8415
rect 14691 8412 14703 8415
rect 15194 8412 15200 8424
rect 14691 8384 15200 8412
rect 14691 8381 14703 8384
rect 14645 8375 14703 8381
rect 15194 8372 15200 8384
rect 15252 8372 15258 8424
rect 15381 8415 15439 8421
rect 15381 8381 15393 8415
rect 15427 8412 15439 8415
rect 16114 8412 16120 8424
rect 15427 8384 16120 8412
rect 15427 8381 15439 8384
rect 15381 8375 15439 8381
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 1104 8186 28888 8208
rect 1104 8134 10243 8186
rect 10295 8134 10307 8186
rect 10359 8134 10371 8186
rect 10423 8134 10435 8186
rect 10487 8134 19504 8186
rect 19556 8134 19568 8186
rect 19620 8134 19632 8186
rect 19684 8134 19696 8186
rect 19748 8134 28888 8186
rect 1104 8112 28888 8134
rect 12342 8072 12348 8084
rect 10796 8044 12348 8072
rect 10796 7945 10824 8044
rect 12342 8032 12348 8044
rect 12400 8072 12406 8084
rect 13265 8075 13323 8081
rect 13265 8072 13277 8075
rect 12400 8044 13277 8072
rect 12400 8032 12406 8044
rect 13265 8041 13277 8044
rect 13311 8041 13323 8075
rect 13265 8035 13323 8041
rect 12158 7964 12164 8016
rect 12216 8004 12222 8016
rect 12621 8007 12679 8013
rect 12621 8004 12633 8007
rect 12216 7976 12633 8004
rect 12216 7964 12222 7976
rect 12621 7973 12633 7976
rect 12667 7973 12679 8007
rect 12621 7967 12679 7973
rect 14734 7964 14740 8016
rect 14792 8004 14798 8016
rect 14982 8007 15040 8013
rect 14982 8004 14994 8007
rect 14792 7976 14994 8004
rect 14792 7964 14798 7976
rect 14982 7973 14994 7976
rect 15028 7973 15040 8007
rect 14982 7967 15040 7973
rect 10781 7939 10839 7945
rect 10781 7905 10793 7939
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7905 11943 7939
rect 12526 7936 12532 7948
rect 12487 7908 12532 7936
rect 11885 7899 11943 7905
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 10594 7868 10600 7880
rect 9824 7840 10600 7868
rect 9824 7828 9830 7840
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 11698 7868 11704 7880
rect 11659 7840 11704 7868
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 11900 7800 11928 7899
rect 12526 7896 12532 7908
rect 12584 7896 12590 7948
rect 12802 7936 12808 7948
rect 12763 7908 12808 7936
rect 12802 7896 12808 7908
rect 12860 7896 12866 7948
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7905 13507 7939
rect 13449 7899 13507 7905
rect 13464 7812 13492 7899
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 14737 7871 14795 7877
rect 14737 7868 14749 7871
rect 13872 7840 14749 7868
rect 13872 7828 13878 7840
rect 14737 7837 14749 7840
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 12250 7800 12256 7812
rect 11900 7772 12256 7800
rect 12250 7760 12256 7772
rect 12308 7800 12314 7812
rect 13446 7800 13452 7812
rect 12308 7772 13452 7800
rect 12308 7760 12314 7772
rect 13446 7760 13452 7772
rect 13504 7760 13510 7812
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 10965 7735 11023 7741
rect 10965 7732 10977 7735
rect 10928 7704 10977 7732
rect 10928 7692 10934 7704
rect 10965 7701 10977 7704
rect 11011 7701 11023 7735
rect 12066 7732 12072 7744
rect 12027 7704 12072 7732
rect 10965 7695 11023 7701
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 12342 7692 12348 7744
rect 12400 7732 12406 7744
rect 12529 7735 12587 7741
rect 12529 7732 12541 7735
rect 12400 7704 12541 7732
rect 12400 7692 12406 7704
rect 12529 7701 12541 7704
rect 12575 7701 12587 7735
rect 12529 7695 12587 7701
rect 15378 7692 15384 7744
rect 15436 7732 15442 7744
rect 16117 7735 16175 7741
rect 16117 7732 16129 7735
rect 15436 7704 16129 7732
rect 15436 7692 15442 7704
rect 16117 7701 16129 7704
rect 16163 7701 16175 7735
rect 16117 7695 16175 7701
rect 1104 7642 28888 7664
rect 1104 7590 5612 7642
rect 5664 7590 5676 7642
rect 5728 7590 5740 7642
rect 5792 7590 5804 7642
rect 5856 7590 14874 7642
rect 14926 7590 14938 7642
rect 14990 7590 15002 7642
rect 15054 7590 15066 7642
rect 15118 7590 24135 7642
rect 24187 7590 24199 7642
rect 24251 7590 24263 7642
rect 24315 7590 24327 7642
rect 24379 7590 28888 7642
rect 1104 7568 28888 7590
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 12250 7528 12256 7540
rect 12211 7500 12256 7528
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 14734 7528 14740 7540
rect 14695 7500 14740 7528
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 15102 7460 15108 7472
rect 14384 7432 15108 7460
rect 13814 7392 13820 7404
rect 12406 7364 13820 7392
rect 10870 7284 10876 7336
rect 10928 7333 10934 7336
rect 10928 7324 10940 7333
rect 10928 7296 10973 7324
rect 10928 7287 10940 7296
rect 10928 7284 10934 7287
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 11112 7296 11161 7324
rect 11112 7284 11118 7296
rect 11149 7293 11161 7296
rect 11195 7324 11207 7327
rect 12406 7324 12434 7364
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 13906 7352 13912 7404
rect 13964 7392 13970 7404
rect 14384 7392 14412 7432
rect 15102 7420 15108 7432
rect 15160 7420 15166 7472
rect 13964 7364 14412 7392
rect 13964 7352 13970 7364
rect 11195 7296 12434 7324
rect 11195 7293 11207 7296
rect 11149 7287 11207 7293
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 14384 7333 14412 7364
rect 15028 7364 15424 7392
rect 14093 7327 14151 7333
rect 14093 7324 14105 7327
rect 13504 7296 14105 7324
rect 13504 7284 13510 7296
rect 14093 7293 14105 7296
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7293 14427 7327
rect 14369 7287 14427 7293
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7324 14519 7327
rect 15028 7324 15056 7364
rect 15396 7336 15424 7364
rect 14507 7296 15056 7324
rect 14507 7293 14519 7296
rect 14461 7287 14519 7293
rect 10594 7216 10600 7268
rect 10652 7256 10658 7268
rect 12069 7259 12127 7265
rect 12069 7256 12081 7259
rect 10652 7228 12081 7256
rect 10652 7216 10658 7228
rect 12069 7225 12081 7228
rect 12115 7225 12127 7259
rect 12069 7219 12127 7225
rect 12285 7259 12343 7265
rect 12285 7225 12297 7259
rect 12331 7256 12343 7259
rect 12894 7256 12900 7268
rect 12331 7228 12900 7256
rect 12331 7225 12343 7228
rect 12285 7219 12343 7225
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 13354 7216 13360 7268
rect 13412 7256 13418 7268
rect 13541 7259 13599 7265
rect 13541 7256 13553 7259
rect 13412 7228 13553 7256
rect 13412 7216 13418 7228
rect 13541 7225 13553 7228
rect 13587 7225 13599 7259
rect 14292 7256 14320 7287
rect 15102 7284 15108 7336
rect 15160 7324 15166 7336
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 15160 7296 15209 7324
rect 15160 7284 15166 7296
rect 15197 7293 15209 7296
rect 15243 7293 15255 7327
rect 15378 7324 15384 7336
rect 15339 7296 15384 7324
rect 15197 7287 15255 7293
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 14550 7256 14556 7268
rect 14292 7228 14556 7256
rect 13541 7219 13599 7225
rect 14550 7216 14556 7228
rect 14608 7256 14614 7268
rect 15289 7259 15347 7265
rect 15289 7256 15301 7259
rect 14608 7228 15301 7256
rect 14608 7216 14614 7228
rect 15289 7225 15301 7228
rect 15335 7225 15347 7259
rect 15289 7219 15347 7225
rect 12437 7191 12495 7197
rect 12437 7157 12449 7191
rect 12483 7188 12495 7191
rect 12710 7188 12716 7200
rect 12483 7160 12716 7188
rect 12483 7157 12495 7160
rect 12437 7151 12495 7157
rect 12710 7148 12716 7160
rect 12768 7148 12774 7200
rect 13449 7191 13507 7197
rect 13449 7157 13461 7191
rect 13495 7188 13507 7191
rect 14458 7188 14464 7200
rect 13495 7160 14464 7188
rect 13495 7157 13507 7160
rect 13449 7151 13507 7157
rect 14458 7148 14464 7160
rect 14516 7188 14522 7200
rect 15010 7188 15016 7200
rect 14516 7160 15016 7188
rect 14516 7148 14522 7160
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 1104 7098 28888 7120
rect 1104 7046 10243 7098
rect 10295 7046 10307 7098
rect 10359 7046 10371 7098
rect 10423 7046 10435 7098
rect 10487 7046 19504 7098
rect 19556 7046 19568 7098
rect 19620 7046 19632 7098
rect 19684 7046 19696 7098
rect 19748 7046 28888 7098
rect 1104 7024 28888 7046
rect 11456 6919 11514 6925
rect 11456 6885 11468 6919
rect 11502 6916 11514 6919
rect 12066 6916 12072 6928
rect 11502 6888 12072 6916
rect 11502 6885 11514 6888
rect 11456 6879 11514 6885
rect 12066 6876 12072 6888
rect 12124 6876 12130 6928
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 10962 6848 10968 6860
rect 10744 6820 10968 6848
rect 10744 6808 10750 6820
rect 10962 6808 10968 6820
rect 11020 6848 11026 6860
rect 11701 6851 11759 6857
rect 11701 6848 11713 6851
rect 11020 6820 11713 6848
rect 11020 6808 11026 6820
rect 11701 6817 11713 6820
rect 11747 6817 11759 6851
rect 11701 6811 11759 6817
rect 12158 6808 12164 6860
rect 12216 6848 12222 6860
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 12216 6820 12265 6848
rect 12216 6808 12222 6820
rect 12253 6817 12265 6820
rect 12299 6817 12311 6851
rect 12253 6811 12311 6817
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 12805 6851 12863 6857
rect 12492 6820 12537 6848
rect 12492 6808 12498 6820
rect 12805 6817 12817 6851
rect 12851 6817 12863 6851
rect 12805 6811 12863 6817
rect 12342 6740 12348 6792
rect 12400 6780 12406 6792
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 12400 6752 12541 6780
rect 12400 6740 12406 6752
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6780 12679 6783
rect 12710 6780 12716 6792
rect 12667 6752 12716 6780
rect 12667 6749 12679 6752
rect 12621 6743 12679 6749
rect 12710 6740 12716 6752
rect 12768 6740 12774 6792
rect 11882 6672 11888 6724
rect 11940 6712 11946 6724
rect 12820 6712 12848 6811
rect 13262 6808 13268 6860
rect 13320 6848 13326 6860
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 13320 6820 13461 6848
rect 13320 6808 13326 6820
rect 13449 6817 13461 6820
rect 13495 6817 13507 6851
rect 13449 6811 13507 6817
rect 13538 6808 13544 6860
rect 13596 6848 13602 6860
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 13596 6820 13645 6848
rect 13596 6808 13602 6820
rect 13633 6817 13645 6820
rect 13679 6817 13691 6851
rect 14921 6851 14979 6857
rect 14921 6848 14933 6851
rect 13633 6811 13691 6817
rect 13740 6820 14933 6848
rect 11940 6684 12848 6712
rect 12989 6715 13047 6721
rect 11940 6672 11946 6684
rect 12544 6656 12572 6684
rect 12989 6681 13001 6715
rect 13035 6712 13047 6715
rect 13630 6712 13636 6724
rect 13035 6684 13636 6712
rect 13035 6681 13047 6684
rect 12989 6675 13047 6681
rect 13630 6672 13636 6684
rect 13688 6672 13694 6724
rect 10321 6647 10379 6653
rect 10321 6613 10333 6647
rect 10367 6644 10379 6647
rect 11054 6644 11060 6656
rect 10367 6616 11060 6644
rect 10367 6613 10379 6616
rect 10321 6607 10379 6613
rect 11054 6604 11060 6616
rect 11112 6644 11118 6656
rect 11698 6644 11704 6656
rect 11112 6616 11704 6644
rect 11112 6604 11118 6616
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 12526 6604 12532 6656
rect 12584 6604 12590 6656
rect 13354 6604 13360 6656
rect 13412 6644 13418 6656
rect 13740 6653 13768 6820
rect 14921 6817 14933 6820
rect 14967 6817 14979 6851
rect 14921 6811 14979 6817
rect 15010 6808 15016 6860
rect 15068 6848 15074 6860
rect 15381 6851 15439 6857
rect 15381 6848 15393 6851
rect 15068 6820 15393 6848
rect 15068 6808 15074 6820
rect 15381 6817 15393 6820
rect 15427 6817 15439 6851
rect 15381 6811 15439 6817
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 14734 6740 14740 6792
rect 14792 6780 14798 6792
rect 15580 6780 15608 6811
rect 14792 6752 15608 6780
rect 14792 6740 14798 6752
rect 13725 6647 13783 6653
rect 13725 6644 13737 6647
rect 13412 6616 13737 6644
rect 13412 6604 13418 6616
rect 13725 6613 13737 6616
rect 13771 6613 13783 6647
rect 13725 6607 13783 6613
rect 14458 6604 14464 6656
rect 14516 6644 14522 6656
rect 14737 6647 14795 6653
rect 14737 6644 14749 6647
rect 14516 6616 14749 6644
rect 14516 6604 14522 6616
rect 14737 6613 14749 6616
rect 14783 6613 14795 6647
rect 15378 6644 15384 6656
rect 15339 6616 15384 6644
rect 14737 6607 14795 6613
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 1104 6554 28888 6576
rect 1104 6502 5612 6554
rect 5664 6502 5676 6554
rect 5728 6502 5740 6554
rect 5792 6502 5804 6554
rect 5856 6502 14874 6554
rect 14926 6502 14938 6554
rect 14990 6502 15002 6554
rect 15054 6502 15066 6554
rect 15118 6502 24135 6554
rect 24187 6502 24199 6554
rect 24251 6502 24263 6554
rect 24315 6502 24327 6554
rect 24379 6502 28888 6554
rect 1104 6480 28888 6502
rect 11149 6443 11207 6449
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11882 6440 11888 6452
rect 11195 6412 11888 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12069 6443 12127 6449
rect 12069 6409 12081 6443
rect 12115 6440 12127 6443
rect 12434 6440 12440 6452
rect 12115 6412 12440 6440
rect 12115 6409 12127 6412
rect 12069 6403 12127 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 13265 6443 13323 6449
rect 13265 6409 13277 6443
rect 13311 6440 13323 6443
rect 13446 6440 13452 6452
rect 13311 6412 13452 6440
rect 13311 6409 13323 6412
rect 13265 6403 13323 6409
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 12636 6276 13952 6304
rect 10134 6236 10140 6248
rect 10095 6208 10140 6236
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 10781 6239 10839 6245
rect 10781 6205 10793 6239
rect 10827 6236 10839 6239
rect 11514 6236 11520 6248
rect 10827 6208 11520 6236
rect 10827 6205 10839 6208
rect 10781 6199 10839 6205
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 12066 6196 12072 6248
rect 12124 6236 12130 6248
rect 12636 6245 12664 6276
rect 12207 6239 12265 6245
rect 12207 6236 12219 6239
rect 12124 6208 12219 6236
rect 12124 6196 12130 6208
rect 12207 6205 12219 6208
rect 12253 6205 12265 6239
rect 12207 6199 12265 6205
rect 12620 6239 12678 6245
rect 12620 6205 12632 6239
rect 12666 6205 12678 6239
rect 12620 6199 12678 6205
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 13354 6236 13360 6248
rect 12768 6208 12813 6236
rect 13315 6208 13360 6236
rect 12768 6196 12774 6208
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 13814 6236 13820 6248
rect 13775 6208 13820 6236
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 13924 6236 13952 6276
rect 14084 6239 14142 6245
rect 14084 6236 14096 6239
rect 13924 6208 14096 6236
rect 14084 6205 14096 6208
rect 14130 6236 14142 6239
rect 15378 6236 15384 6248
rect 14130 6208 15384 6236
rect 14130 6205 14142 6208
rect 14084 6199 14142 6205
rect 15378 6196 15384 6208
rect 15436 6196 15442 6248
rect 10965 6171 11023 6177
rect 10965 6137 10977 6171
rect 11011 6168 11023 6171
rect 11054 6168 11060 6180
rect 11011 6140 11060 6168
rect 11011 6137 11023 6140
rect 10965 6131 11023 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 12342 6168 12348 6180
rect 12303 6140 12348 6168
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 12437 6171 12495 6177
rect 12437 6137 12449 6171
rect 12483 6137 12495 6171
rect 12437 6131 12495 6137
rect 10321 6103 10379 6109
rect 10321 6069 10333 6103
rect 10367 6100 10379 6103
rect 10686 6100 10692 6112
rect 10367 6072 10692 6100
rect 10367 6069 10379 6072
rect 10321 6063 10379 6069
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 12250 6060 12256 6112
rect 12308 6100 12314 6112
rect 12452 6100 12480 6131
rect 13262 6128 13268 6180
rect 13320 6168 13326 6180
rect 16390 6168 16396 6180
rect 13320 6140 16396 6168
rect 13320 6128 13326 6140
rect 16390 6128 16396 6140
rect 16448 6128 16454 6180
rect 12308 6072 12480 6100
rect 12308 6060 12314 6072
rect 14918 6060 14924 6112
rect 14976 6100 14982 6112
rect 15197 6103 15255 6109
rect 15197 6100 15209 6103
rect 14976 6072 15209 6100
rect 14976 6060 14982 6072
rect 15197 6069 15209 6072
rect 15243 6069 15255 6103
rect 15197 6063 15255 6069
rect 1104 6010 28888 6032
rect 1104 5958 10243 6010
rect 10295 5958 10307 6010
rect 10359 5958 10371 6010
rect 10423 5958 10435 6010
rect 10487 5958 19504 6010
rect 19556 5958 19568 6010
rect 19620 5958 19632 6010
rect 19684 5958 19696 6010
rect 19748 5958 28888 6010
rect 1104 5936 28888 5958
rect 11057 5899 11115 5905
rect 11057 5865 11069 5899
rect 11103 5896 11115 5899
rect 12158 5896 12164 5908
rect 11103 5868 12164 5896
rect 11103 5865 11115 5868
rect 11057 5859 11115 5865
rect 12158 5856 12164 5868
rect 12216 5856 12222 5908
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 14734 5896 14740 5908
rect 13872 5868 14740 5896
rect 13872 5856 13878 5868
rect 14734 5856 14740 5868
rect 14792 5896 14798 5908
rect 14829 5899 14887 5905
rect 14829 5896 14841 5899
rect 14792 5868 14841 5896
rect 14792 5856 14798 5868
rect 14829 5865 14841 5868
rect 14875 5865 14887 5899
rect 14829 5859 14887 5865
rect 10594 5788 10600 5840
rect 10652 5828 10658 5840
rect 10873 5831 10931 5837
rect 10873 5828 10885 5831
rect 10652 5800 10885 5828
rect 10652 5788 10658 5800
rect 10873 5797 10885 5800
rect 10919 5797 10931 5831
rect 11514 5828 11520 5840
rect 11475 5800 11520 5828
rect 10873 5791 10931 5797
rect 11514 5788 11520 5800
rect 11572 5788 11578 5840
rect 11701 5831 11759 5837
rect 11701 5797 11713 5831
rect 11747 5828 11759 5831
rect 12342 5828 12348 5840
rect 11747 5800 12348 5828
rect 11747 5797 11759 5800
rect 11701 5791 11759 5797
rect 12342 5788 12348 5800
rect 12400 5788 12406 5840
rect 13354 5828 13360 5840
rect 12544 5800 13360 5828
rect 10689 5763 10747 5769
rect 10689 5729 10701 5763
rect 10735 5729 10747 5763
rect 10689 5723 10747 5729
rect 10042 5652 10048 5704
rect 10100 5692 10106 5704
rect 10704 5692 10732 5723
rect 11146 5720 11152 5772
rect 11204 5760 11210 5772
rect 11885 5763 11943 5769
rect 11885 5760 11897 5763
rect 11204 5732 11897 5760
rect 11204 5720 11210 5732
rect 11885 5729 11897 5732
rect 11931 5760 11943 5763
rect 11974 5760 11980 5772
rect 11931 5732 11980 5760
rect 11931 5729 11943 5732
rect 11885 5723 11943 5729
rect 11974 5720 11980 5732
rect 12032 5760 12038 5772
rect 12544 5769 12572 5800
rect 13354 5788 13360 5800
rect 13412 5788 13418 5840
rect 12529 5763 12587 5769
rect 12032 5732 12480 5760
rect 12032 5720 12038 5732
rect 12345 5695 12403 5701
rect 12345 5692 12357 5695
rect 10100 5664 12357 5692
rect 10100 5652 10106 5664
rect 12345 5661 12357 5664
rect 12391 5661 12403 5695
rect 12345 5655 12403 5661
rect 12452 5624 12480 5732
rect 12529 5729 12541 5763
rect 12575 5729 12587 5763
rect 12529 5723 12587 5729
rect 12713 5763 12771 5769
rect 12713 5729 12725 5763
rect 12759 5760 12771 5763
rect 12894 5760 12900 5772
rect 12759 5732 12900 5760
rect 12759 5729 12771 5732
rect 12713 5723 12771 5729
rect 12894 5720 12900 5732
rect 12952 5720 12958 5772
rect 12986 5720 12992 5772
rect 13044 5760 13050 5772
rect 13265 5763 13323 5769
rect 13265 5760 13277 5763
rect 13044 5732 13277 5760
rect 13044 5720 13050 5732
rect 13265 5729 13277 5732
rect 13311 5729 13323 5763
rect 13265 5723 13323 5729
rect 13449 5763 13507 5769
rect 13449 5729 13461 5763
rect 13495 5760 13507 5763
rect 13906 5760 13912 5772
rect 13495 5732 13912 5760
rect 13495 5729 13507 5732
rect 13449 5723 13507 5729
rect 13906 5720 13912 5732
rect 13964 5720 13970 5772
rect 14918 5760 14924 5772
rect 14879 5732 14924 5760
rect 14918 5720 14924 5732
rect 14976 5720 14982 5772
rect 12912 5692 12940 5720
rect 13633 5695 13691 5701
rect 13633 5692 13645 5695
rect 12912 5664 13645 5692
rect 13633 5661 13645 5664
rect 13679 5661 13691 5695
rect 13633 5655 13691 5661
rect 14458 5624 14464 5636
rect 12452 5596 14464 5624
rect 14458 5584 14464 5596
rect 14516 5584 14522 5636
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 15654 5556 15660 5568
rect 13596 5528 15660 5556
rect 13596 5516 13602 5528
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 1104 5466 28888 5488
rect 1104 5414 5612 5466
rect 5664 5414 5676 5466
rect 5728 5414 5740 5466
rect 5792 5414 5804 5466
rect 5856 5414 14874 5466
rect 14926 5414 14938 5466
rect 14990 5414 15002 5466
rect 15054 5414 15066 5466
rect 15118 5414 24135 5466
rect 24187 5414 24199 5466
rect 24251 5414 24263 5466
rect 24315 5414 24327 5466
rect 24379 5414 28888 5466
rect 1104 5392 28888 5414
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12342 5352 12348 5364
rect 12299 5324 12348 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12802 5312 12808 5364
rect 12860 5352 12866 5364
rect 13265 5355 13323 5361
rect 13265 5352 13277 5355
rect 12860 5324 13277 5352
rect 12860 5312 12866 5324
rect 13265 5321 13277 5324
rect 13311 5321 13323 5355
rect 13265 5315 13323 5321
rect 12268 5256 14320 5284
rect 12268 5228 12296 5256
rect 12250 5176 12256 5228
rect 12308 5176 12314 5228
rect 12526 5216 12532 5228
rect 12487 5188 12532 5216
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 13998 5216 14004 5228
rect 13740 5188 14004 5216
rect 11149 5151 11207 5157
rect 11149 5117 11161 5151
rect 11195 5148 11207 5151
rect 11514 5148 11520 5160
rect 11195 5120 11520 5148
rect 11195 5117 11207 5120
rect 11149 5111 11207 5117
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 12342 5108 12348 5160
rect 12400 5148 12406 5160
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 12400 5120 12449 5148
rect 12400 5108 12406 5120
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 12618 5148 12624 5160
rect 12579 5120 12624 5148
rect 12437 5111 12495 5117
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 12710 5108 12716 5160
rect 12768 5148 12774 5160
rect 13449 5151 13507 5157
rect 12768 5120 12813 5148
rect 12768 5108 12774 5120
rect 13449 5117 13461 5151
rect 13495 5117 13507 5151
rect 13449 5111 13507 5117
rect 13541 5151 13599 5157
rect 13541 5117 13553 5151
rect 13587 5148 13599 5151
rect 13630 5148 13636 5160
rect 13587 5120 13636 5148
rect 13587 5117 13599 5120
rect 13541 5111 13599 5117
rect 13464 5080 13492 5111
rect 13630 5108 13636 5120
rect 13688 5108 13694 5160
rect 13740 5157 13768 5188
rect 13998 5176 14004 5188
rect 14056 5176 14062 5228
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5117 13783 5151
rect 13725 5111 13783 5117
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 14292 5157 14320 5256
rect 14277 5151 14335 5157
rect 13872 5120 13917 5148
rect 13872 5108 13878 5120
rect 14277 5117 14289 5151
rect 14323 5117 14335 5151
rect 14458 5148 14464 5160
rect 14419 5120 14464 5148
rect 14277 5111 14335 5117
rect 14458 5108 14464 5120
rect 14516 5108 14522 5160
rect 15930 5148 15936 5160
rect 15891 5120 15936 5148
rect 15930 5108 15936 5120
rect 15988 5108 15994 5160
rect 14369 5083 14427 5089
rect 14369 5080 14381 5083
rect 13464 5052 14381 5080
rect 13556 5024 13584 5052
rect 14369 5049 14381 5052
rect 14415 5049 14427 5083
rect 14369 5043 14427 5049
rect 11054 5012 11060 5024
rect 11015 4984 11060 5012
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 13538 4972 13544 5024
rect 13596 4972 13602 5024
rect 15841 5015 15899 5021
rect 15841 4981 15853 5015
rect 15887 5012 15899 5015
rect 16206 5012 16212 5024
rect 15887 4984 16212 5012
rect 15887 4981 15899 4984
rect 15841 4975 15899 4981
rect 16206 4972 16212 4984
rect 16264 4972 16270 5024
rect 1104 4922 28888 4944
rect 1104 4870 10243 4922
rect 10295 4870 10307 4922
rect 10359 4870 10371 4922
rect 10423 4870 10435 4922
rect 10487 4870 19504 4922
rect 19556 4870 19568 4922
rect 19620 4870 19632 4922
rect 19684 4870 19696 4922
rect 19748 4870 28888 4922
rect 1104 4848 28888 4870
rect 12710 4817 12716 4820
rect 11885 4811 11943 4817
rect 11885 4777 11897 4811
rect 11931 4777 11943 4811
rect 12706 4808 12716 4817
rect 12671 4780 12716 4808
rect 11885 4771 11943 4777
rect 12706 4771 12716 4780
rect 10772 4743 10830 4749
rect 10772 4709 10784 4743
rect 10818 4740 10830 4743
rect 11054 4740 11060 4752
rect 10818 4712 11060 4740
rect 10818 4709 10830 4712
rect 10772 4703 10830 4709
rect 11054 4700 11060 4712
rect 11112 4700 11118 4752
rect 11900 4740 11928 4771
rect 12710 4768 12716 4771
rect 12768 4768 12774 4820
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 13541 4811 13599 4817
rect 13541 4808 13553 4811
rect 12952 4780 13553 4808
rect 12952 4768 12958 4780
rect 13541 4777 13553 4780
rect 13587 4777 13599 4811
rect 13541 4771 13599 4777
rect 13817 4811 13875 4817
rect 13817 4777 13829 4811
rect 13863 4808 13875 4811
rect 13906 4808 13912 4820
rect 13863 4780 13912 4808
rect 13863 4777 13875 4780
rect 13817 4771 13875 4777
rect 13906 4768 13912 4780
rect 13964 4768 13970 4820
rect 16206 4808 16212 4820
rect 16167 4780 16212 4808
rect 16206 4768 16212 4780
rect 16264 4768 16270 4820
rect 12158 4740 12164 4752
rect 11900 4712 12164 4740
rect 12158 4700 12164 4712
rect 12216 4740 12222 4752
rect 12342 4740 12348 4752
rect 12216 4712 12348 4740
rect 12216 4700 12222 4712
rect 12342 4700 12348 4712
rect 12400 4740 12406 4752
rect 12805 4743 12863 4749
rect 12805 4740 12817 4743
rect 12400 4712 12817 4740
rect 12400 4700 12406 4712
rect 12805 4709 12817 4712
rect 12851 4740 12863 4743
rect 13633 4743 13691 4749
rect 13633 4740 13645 4743
rect 12851 4712 13645 4740
rect 12851 4709 12863 4712
rect 12805 4703 12863 4709
rect 13633 4709 13645 4712
rect 13679 4709 13691 4743
rect 13633 4703 13691 4709
rect 10042 4672 10048 4684
rect 10003 4644 10048 4672
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 10505 4675 10563 4681
rect 10505 4641 10517 4675
rect 10551 4672 10563 4675
rect 10594 4672 10600 4684
rect 10551 4644 10600 4672
rect 10551 4641 10563 4644
rect 10505 4635 10563 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 12526 4672 12532 4684
rect 12487 4644 12532 4672
rect 12526 4632 12532 4644
rect 12584 4632 12590 4684
rect 12618 4632 12624 4684
rect 12676 4672 12682 4684
rect 13449 4675 13507 4681
rect 12676 4644 12721 4672
rect 12676 4632 12682 4644
rect 13449 4641 13461 4675
rect 13495 4641 13507 4675
rect 13449 4635 13507 4641
rect 12342 4564 12348 4616
rect 12400 4604 12406 4616
rect 13464 4604 13492 4635
rect 13998 4632 14004 4684
rect 14056 4672 14062 4684
rect 14734 4672 14740 4684
rect 14056 4644 14740 4672
rect 14056 4632 14062 4644
rect 14734 4632 14740 4644
rect 14792 4632 14798 4684
rect 16301 4675 16359 4681
rect 16301 4641 16313 4675
rect 16347 4672 16359 4675
rect 17862 4672 17868 4684
rect 16347 4644 17868 4672
rect 16347 4641 16359 4644
rect 16301 4635 16359 4641
rect 17862 4632 17868 4644
rect 17920 4632 17926 4684
rect 14366 4604 14372 4616
rect 12400 4576 14372 4604
rect 12400 4564 12406 4576
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 16390 4604 16396 4616
rect 16351 4576 16396 4604
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 13262 4536 13268 4548
rect 13223 4508 13268 4536
rect 13262 4496 13268 4508
rect 13320 4496 13326 4548
rect 9950 4468 9956 4480
rect 9911 4440 9956 4468
rect 9950 4428 9956 4440
rect 10008 4428 10014 4480
rect 14829 4471 14887 4477
rect 14829 4437 14841 4471
rect 14875 4468 14887 4471
rect 15286 4468 15292 4480
rect 14875 4440 15292 4468
rect 14875 4437 14887 4440
rect 14829 4431 14887 4437
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 15838 4468 15844 4480
rect 15799 4440 15844 4468
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 1104 4378 28888 4400
rect 1104 4326 5612 4378
rect 5664 4326 5676 4378
rect 5728 4326 5740 4378
rect 5792 4326 5804 4378
rect 5856 4326 14874 4378
rect 14926 4326 14938 4378
rect 14990 4326 15002 4378
rect 15054 4326 15066 4378
rect 15118 4326 24135 4378
rect 24187 4326 24199 4378
rect 24251 4326 24263 4378
rect 24315 4326 24327 4378
rect 24379 4326 28888 4378
rect 1104 4304 28888 4326
rect 12526 4264 12532 4276
rect 12084 4236 12532 4264
rect 12084 4128 12112 4236
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 14366 4264 14372 4276
rect 14327 4236 14372 4264
rect 14366 4224 14372 4236
rect 14424 4224 14430 4276
rect 15930 4224 15936 4276
rect 15988 4264 15994 4276
rect 16393 4267 16451 4273
rect 16393 4264 16405 4267
rect 15988 4236 16405 4264
rect 15988 4224 15994 4236
rect 16393 4233 16405 4236
rect 16439 4233 16451 4267
rect 16393 4227 16451 4233
rect 12802 4196 12808 4208
rect 10980 4100 12112 4128
rect 12268 4168 12808 4196
rect 10980 4069 11008 4100
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4029 11023 4063
rect 11146 4060 11152 4072
rect 11107 4032 11152 4060
rect 10965 4023 11023 4029
rect 11146 4020 11152 4032
rect 11204 4020 11210 4072
rect 12158 4060 12164 4072
rect 12119 4032 12164 4060
rect 12158 4020 12164 4032
rect 12216 4020 12222 4072
rect 10594 3952 10600 4004
rect 10652 3992 10658 4004
rect 11790 3992 11796 4004
rect 10652 3964 11796 3992
rect 10652 3952 10658 3964
rect 11790 3952 11796 3964
rect 11848 3952 11854 4004
rect 12268 3992 12296 4168
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 12387 4131 12445 4137
rect 12387 4097 12399 4131
rect 12433 4128 12445 4131
rect 12618 4128 12624 4140
rect 12433 4100 12624 4128
rect 12433 4097 12445 4100
rect 12387 4091 12445 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4060 12587 4063
rect 12894 4060 12900 4072
rect 12575 4032 12900 4060
rect 12575 4029 12587 4032
rect 12529 4023 12587 4029
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 12989 4063 13047 4069
rect 12989 4029 13001 4063
rect 13035 4060 13047 4063
rect 13814 4060 13820 4072
rect 13035 4032 13820 4060
rect 13035 4029 13047 4032
rect 12989 4023 13047 4029
rect 13814 4020 13820 4032
rect 13872 4060 13878 4072
rect 15286 4069 15292 4072
rect 15013 4063 15071 4069
rect 15013 4060 15025 4063
rect 13872 4032 15025 4060
rect 13872 4020 13878 4032
rect 15013 4029 15025 4032
rect 15059 4029 15071 4063
rect 15280 4060 15292 4069
rect 15247 4032 15292 4060
rect 15013 4023 15071 4029
rect 15280 4023 15292 4032
rect 15286 4020 15292 4023
rect 15344 4020 15350 4072
rect 12176 3964 12296 3992
rect 11057 3927 11115 3933
rect 11057 3893 11069 3927
rect 11103 3924 11115 3927
rect 12176 3924 12204 3964
rect 12802 3952 12808 4004
rect 12860 3992 12866 4004
rect 13234 3995 13292 4001
rect 13234 3992 13246 3995
rect 12860 3964 13246 3992
rect 12860 3952 12866 3964
rect 13234 3961 13246 3964
rect 13280 3992 13292 3995
rect 13722 3992 13728 4004
rect 13280 3964 13728 3992
rect 13280 3961 13292 3964
rect 13234 3955 13292 3961
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 11103 3896 12204 3924
rect 12253 3927 12311 3933
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 12253 3893 12265 3927
rect 12299 3924 12311 3927
rect 12342 3924 12348 3936
rect 12299 3896 12348 3924
rect 12299 3893 12311 3896
rect 12253 3887 12311 3893
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 12986 3924 12992 3936
rect 12483 3896 12992 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 1104 3834 28888 3856
rect 1104 3782 10243 3834
rect 10295 3782 10307 3834
rect 10359 3782 10371 3834
rect 10423 3782 10435 3834
rect 10487 3782 19504 3834
rect 19556 3782 19568 3834
rect 19620 3782 19632 3834
rect 19684 3782 19696 3834
rect 19748 3782 28888 3834
rect 1104 3760 28888 3782
rect 12437 3723 12495 3729
rect 12437 3689 12449 3723
rect 12483 3720 12495 3723
rect 13262 3720 13268 3732
rect 12483 3692 13268 3720
rect 12483 3689 12495 3692
rect 12437 3683 12495 3689
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 15105 3723 15163 3729
rect 15105 3720 15117 3723
rect 14792 3692 15117 3720
rect 14792 3680 14798 3692
rect 15105 3689 15117 3692
rect 15151 3689 15163 3723
rect 15105 3683 15163 3689
rect 15473 3723 15531 3729
rect 15473 3689 15485 3723
rect 15519 3720 15531 3723
rect 15838 3720 15844 3732
rect 15519 3692 15844 3720
rect 15519 3689 15531 3692
rect 15473 3683 15531 3689
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 10842 3655 10900 3661
rect 10842 3652 10854 3655
rect 10008 3624 10854 3652
rect 10008 3612 10014 3624
rect 10842 3621 10854 3624
rect 10888 3621 10900 3655
rect 10842 3615 10900 3621
rect 12406 3624 13860 3652
rect 10597 3587 10655 3593
rect 10597 3553 10609 3587
rect 10643 3584 10655 3587
rect 10686 3584 10692 3596
rect 10643 3556 10692 3584
rect 10643 3553 10655 3556
rect 10597 3547 10655 3553
rect 10686 3544 10692 3556
rect 10744 3584 10750 3596
rect 12406 3584 12434 3624
rect 13832 3596 13860 3624
rect 10744 3556 12434 3584
rect 10744 3544 10750 3556
rect 13538 3544 13544 3596
rect 13596 3593 13602 3596
rect 13596 3584 13608 3593
rect 13814 3584 13820 3596
rect 13596 3556 13641 3584
rect 13775 3556 13820 3584
rect 13596 3547 13608 3556
rect 13596 3544 13602 3547
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 15565 3587 15623 3593
rect 15565 3553 15577 3587
rect 15611 3584 15623 3587
rect 15611 3556 22094 3584
rect 15611 3553 15623 3556
rect 15565 3547 15623 3553
rect 15654 3516 15660 3528
rect 15615 3488 15660 3516
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 22066 3516 22094 3556
rect 27890 3516 27896 3528
rect 22066 3488 27896 3516
rect 27890 3476 27896 3488
rect 27948 3476 27954 3528
rect 11977 3383 12035 3389
rect 11977 3349 11989 3383
rect 12023 3380 12035 3383
rect 12894 3380 12900 3392
rect 12023 3352 12900 3380
rect 12023 3349 12035 3352
rect 11977 3343 12035 3349
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 1104 3290 28888 3312
rect 1104 3238 5612 3290
rect 5664 3238 5676 3290
rect 5728 3238 5740 3290
rect 5792 3238 5804 3290
rect 5856 3238 14874 3290
rect 14926 3238 14938 3290
rect 14990 3238 15002 3290
rect 15054 3238 15066 3290
rect 15118 3238 24135 3290
rect 24187 3238 24199 3290
rect 24251 3238 24263 3290
rect 24315 3238 24327 3290
rect 24379 3238 28888 3290
rect 1104 3216 28888 3238
rect 12250 3136 12256 3188
rect 12308 3176 12314 3188
rect 12345 3179 12403 3185
rect 12345 3176 12357 3179
rect 12308 3148 12357 3176
rect 12308 3136 12314 3148
rect 12345 3145 12357 3148
rect 12391 3145 12403 3179
rect 12345 3139 12403 3145
rect 17862 3136 17868 3188
rect 17920 3176 17926 3188
rect 19889 3179 19947 3185
rect 19889 3176 19901 3179
rect 17920 3148 19901 3176
rect 17920 3136 17926 3148
rect 19889 3145 19901 3148
rect 19935 3145 19947 3179
rect 27890 3176 27896 3188
rect 27851 3148 27896 3176
rect 19889 3139 19947 3145
rect 27890 3136 27896 3148
rect 27948 3136 27954 3188
rect 13173 3111 13231 3117
rect 13173 3077 13185 3111
rect 13219 3108 13231 3111
rect 13909 3111 13967 3117
rect 13909 3108 13921 3111
rect 13219 3080 13921 3108
rect 13219 3077 13231 3080
rect 13173 3071 13231 3077
rect 13909 3077 13921 3080
rect 13955 3077 13967 3111
rect 13909 3071 13967 3077
rect 12618 3040 12624 3052
rect 12176 3012 12624 3040
rect 12176 2981 12204 3012
rect 12618 3000 12624 3012
rect 12676 3040 12682 3052
rect 12676 3012 12756 3040
rect 12676 3000 12682 3012
rect 12161 2975 12219 2981
rect 12161 2941 12173 2975
rect 12207 2941 12219 2975
rect 12161 2935 12219 2941
rect 12345 2975 12403 2981
rect 12345 2941 12357 2975
rect 12391 2972 12403 2975
rect 12526 2972 12532 2984
rect 12391 2944 12532 2972
rect 12391 2941 12403 2944
rect 12345 2935 12403 2941
rect 12526 2932 12532 2944
rect 12584 2972 12590 2984
rect 12728 2981 12756 3012
rect 12713 2975 12771 2981
rect 12584 2944 12664 2972
rect 12584 2932 12590 2944
rect 12636 2845 12664 2944
rect 12713 2941 12725 2975
rect 12759 2941 12771 2975
rect 12713 2935 12771 2941
rect 12728 2904 12756 2935
rect 13262 2932 13268 2984
rect 13320 2972 13326 2984
rect 13449 2975 13507 2981
rect 13449 2972 13461 2975
rect 13320 2944 13461 2972
rect 13320 2932 13326 2944
rect 13449 2941 13461 2944
rect 13495 2941 13507 2975
rect 13449 2935 13507 2941
rect 14093 2975 14151 2981
rect 14093 2941 14105 2975
rect 14139 2972 14151 2975
rect 14366 2972 14372 2984
rect 14139 2944 14372 2972
rect 14139 2941 14151 2944
rect 14093 2935 14151 2941
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 19981 2975 20039 2981
rect 19981 2941 19993 2975
rect 20027 2972 20039 2975
rect 20714 2972 20720 2984
rect 20027 2944 20720 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 20714 2932 20720 2944
rect 20772 2932 20778 2984
rect 27338 2932 27344 2984
rect 27396 2972 27402 2984
rect 27801 2975 27859 2981
rect 27801 2972 27813 2975
rect 27396 2944 27813 2972
rect 27396 2932 27402 2944
rect 27801 2941 27813 2944
rect 27847 2941 27859 2975
rect 27801 2935 27859 2941
rect 12728 2876 13308 2904
rect 13280 2845 13308 2876
rect 12621 2839 12679 2845
rect 12621 2805 12633 2839
rect 12667 2836 12679 2839
rect 13173 2839 13231 2845
rect 13173 2836 13185 2839
rect 12667 2808 13185 2836
rect 12667 2805 12679 2808
rect 12621 2799 12679 2805
rect 13173 2805 13185 2808
rect 13219 2805 13231 2839
rect 13173 2799 13231 2805
rect 13265 2839 13323 2845
rect 13265 2805 13277 2839
rect 13311 2805 13323 2839
rect 13265 2799 13323 2805
rect 1104 2746 28888 2768
rect 1104 2694 10243 2746
rect 10295 2694 10307 2746
rect 10359 2694 10371 2746
rect 10423 2694 10435 2746
rect 10487 2694 19504 2746
rect 19556 2694 19568 2746
rect 19620 2694 19632 2746
rect 19684 2694 19696 2746
rect 19748 2694 28888 2746
rect 1104 2672 28888 2694
rect 1578 2632 1584 2644
rect 1539 2604 1584 2632
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 20714 2632 20720 2644
rect 20675 2604 20720 2632
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 27338 2632 27344 2644
rect 27299 2604 27344 2632
rect 27338 2592 27344 2604
rect 27396 2592 27402 2644
rect 474 2456 480 2508
rect 532 2496 538 2508
rect 1397 2499 1455 2505
rect 1397 2496 1409 2499
rect 532 2468 1409 2496
rect 532 2456 538 2468
rect 1397 2465 1409 2468
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 20714 2456 20720 2508
rect 20772 2496 20778 2508
rect 20901 2499 20959 2505
rect 20901 2496 20913 2499
rect 20772 2468 20913 2496
rect 20772 2456 20778 2468
rect 20901 2465 20913 2468
rect 20947 2465 20959 2499
rect 27154 2496 27160 2508
rect 27115 2468 27160 2496
rect 20901 2459 20959 2465
rect 27154 2456 27160 2468
rect 27212 2456 27218 2508
rect 1104 2202 28888 2224
rect 1104 2150 5612 2202
rect 5664 2150 5676 2202
rect 5728 2150 5740 2202
rect 5792 2150 5804 2202
rect 5856 2150 14874 2202
rect 14926 2150 14938 2202
rect 14990 2150 15002 2202
rect 15054 2150 15066 2202
rect 15118 2150 24135 2202
rect 24187 2150 24199 2202
rect 24251 2150 24263 2202
rect 24315 2150 24327 2202
rect 24379 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 10243 29894 10295 29946
rect 10307 29894 10359 29946
rect 10371 29894 10423 29946
rect 10435 29894 10487 29946
rect 19504 29894 19556 29946
rect 19568 29894 19620 29946
rect 19632 29894 19684 29946
rect 19696 29894 19748 29946
rect 29460 29724 29512 29776
rect 1400 29699 1452 29708
rect 1400 29665 1409 29699
rect 1409 29665 1443 29699
rect 1443 29665 1452 29699
rect 1400 29656 1452 29665
rect 9220 29656 9272 29708
rect 19340 29699 19392 29708
rect 19340 29665 19349 29699
rect 19349 29665 19383 29699
rect 19383 29665 19392 29699
rect 19340 29656 19392 29665
rect 1584 29495 1636 29504
rect 1584 29461 1593 29495
rect 1593 29461 1627 29495
rect 1627 29461 1636 29495
rect 1584 29452 1636 29461
rect 9772 29495 9824 29504
rect 9772 29461 9781 29495
rect 9781 29461 9815 29495
rect 9815 29461 9824 29495
rect 9772 29452 9824 29461
rect 14740 29452 14792 29504
rect 5612 29350 5664 29402
rect 5676 29350 5728 29402
rect 5740 29350 5792 29402
rect 5804 29350 5856 29402
rect 14874 29350 14926 29402
rect 14938 29350 14990 29402
rect 15002 29350 15054 29402
rect 15066 29350 15118 29402
rect 24135 29350 24187 29402
rect 24199 29350 24251 29402
rect 24263 29350 24315 29402
rect 24327 29350 24379 29402
rect 10243 28806 10295 28858
rect 10307 28806 10359 28858
rect 10371 28806 10423 28858
rect 10435 28806 10487 28858
rect 19504 28806 19556 28858
rect 19568 28806 19620 28858
rect 19632 28806 19684 28858
rect 19696 28806 19748 28858
rect 5612 28262 5664 28314
rect 5676 28262 5728 28314
rect 5740 28262 5792 28314
rect 5804 28262 5856 28314
rect 14874 28262 14926 28314
rect 14938 28262 14990 28314
rect 15002 28262 15054 28314
rect 15066 28262 15118 28314
rect 24135 28262 24187 28314
rect 24199 28262 24251 28314
rect 24263 28262 24315 28314
rect 24327 28262 24379 28314
rect 10243 27718 10295 27770
rect 10307 27718 10359 27770
rect 10371 27718 10423 27770
rect 10435 27718 10487 27770
rect 19504 27718 19556 27770
rect 19568 27718 19620 27770
rect 19632 27718 19684 27770
rect 19696 27718 19748 27770
rect 5612 27174 5664 27226
rect 5676 27174 5728 27226
rect 5740 27174 5792 27226
rect 5804 27174 5856 27226
rect 14874 27174 14926 27226
rect 14938 27174 14990 27226
rect 15002 27174 15054 27226
rect 15066 27174 15118 27226
rect 24135 27174 24187 27226
rect 24199 27174 24251 27226
rect 24263 27174 24315 27226
rect 24327 27174 24379 27226
rect 10243 26630 10295 26682
rect 10307 26630 10359 26682
rect 10371 26630 10423 26682
rect 10435 26630 10487 26682
rect 19504 26630 19556 26682
rect 19568 26630 19620 26682
rect 19632 26630 19684 26682
rect 19696 26630 19748 26682
rect 5612 26086 5664 26138
rect 5676 26086 5728 26138
rect 5740 26086 5792 26138
rect 5804 26086 5856 26138
rect 14874 26086 14926 26138
rect 14938 26086 14990 26138
rect 15002 26086 15054 26138
rect 15066 26086 15118 26138
rect 24135 26086 24187 26138
rect 24199 26086 24251 26138
rect 24263 26086 24315 26138
rect 24327 26086 24379 26138
rect 10243 25542 10295 25594
rect 10307 25542 10359 25594
rect 10371 25542 10423 25594
rect 10435 25542 10487 25594
rect 19504 25542 19556 25594
rect 19568 25542 19620 25594
rect 19632 25542 19684 25594
rect 19696 25542 19748 25594
rect 5612 24998 5664 25050
rect 5676 24998 5728 25050
rect 5740 24998 5792 25050
rect 5804 24998 5856 25050
rect 14874 24998 14926 25050
rect 14938 24998 14990 25050
rect 15002 24998 15054 25050
rect 15066 24998 15118 25050
rect 24135 24998 24187 25050
rect 24199 24998 24251 25050
rect 24263 24998 24315 25050
rect 24327 24998 24379 25050
rect 10243 24454 10295 24506
rect 10307 24454 10359 24506
rect 10371 24454 10423 24506
rect 10435 24454 10487 24506
rect 19504 24454 19556 24506
rect 19568 24454 19620 24506
rect 19632 24454 19684 24506
rect 19696 24454 19748 24506
rect 5612 23910 5664 23962
rect 5676 23910 5728 23962
rect 5740 23910 5792 23962
rect 5804 23910 5856 23962
rect 14874 23910 14926 23962
rect 14938 23910 14990 23962
rect 15002 23910 15054 23962
rect 15066 23910 15118 23962
rect 24135 23910 24187 23962
rect 24199 23910 24251 23962
rect 24263 23910 24315 23962
rect 24327 23910 24379 23962
rect 10243 23366 10295 23418
rect 10307 23366 10359 23418
rect 10371 23366 10423 23418
rect 10435 23366 10487 23418
rect 19504 23366 19556 23418
rect 19568 23366 19620 23418
rect 19632 23366 19684 23418
rect 19696 23366 19748 23418
rect 5612 22822 5664 22874
rect 5676 22822 5728 22874
rect 5740 22822 5792 22874
rect 5804 22822 5856 22874
rect 14874 22822 14926 22874
rect 14938 22822 14990 22874
rect 15002 22822 15054 22874
rect 15066 22822 15118 22874
rect 24135 22822 24187 22874
rect 24199 22822 24251 22874
rect 24263 22822 24315 22874
rect 24327 22822 24379 22874
rect 10243 22278 10295 22330
rect 10307 22278 10359 22330
rect 10371 22278 10423 22330
rect 10435 22278 10487 22330
rect 19504 22278 19556 22330
rect 19568 22278 19620 22330
rect 19632 22278 19684 22330
rect 19696 22278 19748 22330
rect 5612 21734 5664 21786
rect 5676 21734 5728 21786
rect 5740 21734 5792 21786
rect 5804 21734 5856 21786
rect 14874 21734 14926 21786
rect 14938 21734 14990 21786
rect 15002 21734 15054 21786
rect 15066 21734 15118 21786
rect 24135 21734 24187 21786
rect 24199 21734 24251 21786
rect 24263 21734 24315 21786
rect 24327 21734 24379 21786
rect 10243 21190 10295 21242
rect 10307 21190 10359 21242
rect 10371 21190 10423 21242
rect 10435 21190 10487 21242
rect 19504 21190 19556 21242
rect 19568 21190 19620 21242
rect 19632 21190 19684 21242
rect 19696 21190 19748 21242
rect 5612 20646 5664 20698
rect 5676 20646 5728 20698
rect 5740 20646 5792 20698
rect 5804 20646 5856 20698
rect 14874 20646 14926 20698
rect 14938 20646 14990 20698
rect 15002 20646 15054 20698
rect 15066 20646 15118 20698
rect 24135 20646 24187 20698
rect 24199 20646 24251 20698
rect 24263 20646 24315 20698
rect 24327 20646 24379 20698
rect 10243 20102 10295 20154
rect 10307 20102 10359 20154
rect 10371 20102 10423 20154
rect 10435 20102 10487 20154
rect 19504 20102 19556 20154
rect 19568 20102 19620 20154
rect 19632 20102 19684 20154
rect 19696 20102 19748 20154
rect 5612 19558 5664 19610
rect 5676 19558 5728 19610
rect 5740 19558 5792 19610
rect 5804 19558 5856 19610
rect 14874 19558 14926 19610
rect 14938 19558 14990 19610
rect 15002 19558 15054 19610
rect 15066 19558 15118 19610
rect 24135 19558 24187 19610
rect 24199 19558 24251 19610
rect 24263 19558 24315 19610
rect 24327 19558 24379 19610
rect 10243 19014 10295 19066
rect 10307 19014 10359 19066
rect 10371 19014 10423 19066
rect 10435 19014 10487 19066
rect 19504 19014 19556 19066
rect 19568 19014 19620 19066
rect 19632 19014 19684 19066
rect 19696 19014 19748 19066
rect 5612 18470 5664 18522
rect 5676 18470 5728 18522
rect 5740 18470 5792 18522
rect 5804 18470 5856 18522
rect 14874 18470 14926 18522
rect 14938 18470 14990 18522
rect 15002 18470 15054 18522
rect 15066 18470 15118 18522
rect 24135 18470 24187 18522
rect 24199 18470 24251 18522
rect 24263 18470 24315 18522
rect 24327 18470 24379 18522
rect 10243 17926 10295 17978
rect 10307 17926 10359 17978
rect 10371 17926 10423 17978
rect 10435 17926 10487 17978
rect 19504 17926 19556 17978
rect 19568 17926 19620 17978
rect 19632 17926 19684 17978
rect 19696 17926 19748 17978
rect 5612 17382 5664 17434
rect 5676 17382 5728 17434
rect 5740 17382 5792 17434
rect 5804 17382 5856 17434
rect 14874 17382 14926 17434
rect 14938 17382 14990 17434
rect 15002 17382 15054 17434
rect 15066 17382 15118 17434
rect 24135 17382 24187 17434
rect 24199 17382 24251 17434
rect 24263 17382 24315 17434
rect 24327 17382 24379 17434
rect 27988 17051 28040 17060
rect 27988 17017 27997 17051
rect 27997 17017 28031 17051
rect 28031 17017 28040 17051
rect 27988 17008 28040 17017
rect 28172 17051 28224 17060
rect 28172 17017 28181 17051
rect 28181 17017 28215 17051
rect 28215 17017 28224 17051
rect 28172 17008 28224 17017
rect 10243 16838 10295 16890
rect 10307 16838 10359 16890
rect 10371 16838 10423 16890
rect 10435 16838 10487 16890
rect 19504 16838 19556 16890
rect 19568 16838 19620 16890
rect 19632 16838 19684 16890
rect 19696 16838 19748 16890
rect 5612 16294 5664 16346
rect 5676 16294 5728 16346
rect 5740 16294 5792 16346
rect 5804 16294 5856 16346
rect 14874 16294 14926 16346
rect 14938 16294 14990 16346
rect 15002 16294 15054 16346
rect 15066 16294 15118 16346
rect 24135 16294 24187 16346
rect 24199 16294 24251 16346
rect 24263 16294 24315 16346
rect 24327 16294 24379 16346
rect 10243 15750 10295 15802
rect 10307 15750 10359 15802
rect 10371 15750 10423 15802
rect 10435 15750 10487 15802
rect 19504 15750 19556 15802
rect 19568 15750 19620 15802
rect 19632 15750 19684 15802
rect 19696 15750 19748 15802
rect 14740 15512 14792 15564
rect 13820 15308 13872 15360
rect 5612 15206 5664 15258
rect 5676 15206 5728 15258
rect 5740 15206 5792 15258
rect 5804 15206 5856 15258
rect 14874 15206 14926 15258
rect 14938 15206 14990 15258
rect 15002 15206 15054 15258
rect 15066 15206 15118 15258
rect 24135 15206 24187 15258
rect 24199 15206 24251 15258
rect 24263 15206 24315 15258
rect 24327 15206 24379 15258
rect 1584 14968 1636 15020
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 12256 14900 12308 14952
rect 12900 14900 12952 14952
rect 8484 14764 8536 14816
rect 12808 14764 12860 14816
rect 13820 14900 13872 14952
rect 13728 14764 13780 14816
rect 10243 14662 10295 14714
rect 10307 14662 10359 14714
rect 10371 14662 10423 14714
rect 10435 14662 10487 14714
rect 19504 14662 19556 14714
rect 19568 14662 19620 14714
rect 19632 14662 19684 14714
rect 19696 14662 19748 14714
rect 8484 14492 8536 14544
rect 12256 14424 12308 14476
rect 12808 14467 12860 14476
rect 12808 14433 12817 14467
rect 12817 14433 12851 14467
rect 12851 14433 12860 14467
rect 12808 14424 12860 14433
rect 13820 14424 13872 14476
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 13084 14288 13136 14340
rect 13544 14220 13596 14272
rect 5612 14118 5664 14170
rect 5676 14118 5728 14170
rect 5740 14118 5792 14170
rect 5804 14118 5856 14170
rect 14874 14118 14926 14170
rect 14938 14118 14990 14170
rect 15002 14118 15054 14170
rect 15066 14118 15118 14170
rect 24135 14118 24187 14170
rect 24199 14118 24251 14170
rect 24263 14118 24315 14170
rect 24327 14118 24379 14170
rect 12072 13948 12124 14000
rect 13176 13855 13228 13864
rect 13176 13821 13194 13855
rect 13194 13821 13228 13855
rect 13176 13812 13228 13821
rect 13452 13855 13504 13864
rect 13452 13821 13461 13855
rect 13461 13821 13495 13855
rect 13495 13821 13504 13855
rect 13452 13812 13504 13821
rect 12900 13744 12952 13796
rect 14372 13744 14424 13796
rect 12164 13676 12216 13728
rect 15292 13719 15344 13728
rect 15292 13685 15301 13719
rect 15301 13685 15335 13719
rect 15335 13685 15344 13719
rect 27988 13812 28040 13864
rect 15292 13676 15344 13685
rect 10243 13574 10295 13626
rect 10307 13574 10359 13626
rect 10371 13574 10423 13626
rect 10435 13574 10487 13626
rect 19504 13574 19556 13626
rect 19568 13574 19620 13626
rect 19632 13574 19684 13626
rect 19696 13574 19748 13626
rect 12256 13472 12308 13524
rect 1584 13336 1636 13388
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 12900 13336 12952 13388
rect 15292 13336 15344 13388
rect 9772 13268 9824 13320
rect 12072 13311 12124 13320
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 13084 13268 13136 13320
rect 14004 13132 14056 13184
rect 5612 13030 5664 13082
rect 5676 13030 5728 13082
rect 5740 13030 5792 13082
rect 5804 13030 5856 13082
rect 14874 13030 14926 13082
rect 14938 13030 14990 13082
rect 15002 13030 15054 13082
rect 15066 13030 15118 13082
rect 24135 13030 24187 13082
rect 24199 13030 24251 13082
rect 24263 13030 24315 13082
rect 24327 13030 24379 13082
rect 13084 12928 13136 12980
rect 14372 12971 14424 12980
rect 14372 12937 14381 12971
rect 14381 12937 14415 12971
rect 14415 12937 14424 12971
rect 14372 12928 14424 12937
rect 9956 12724 10008 12776
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 12164 12767 12216 12776
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 14004 12767 14056 12776
rect 14004 12733 14013 12767
rect 14013 12733 14047 12767
rect 14047 12733 14056 12767
rect 14004 12724 14056 12733
rect 12624 12656 12676 12708
rect 14556 12656 14608 12708
rect 12532 12588 12584 12640
rect 10243 12486 10295 12538
rect 10307 12486 10359 12538
rect 10371 12486 10423 12538
rect 10435 12486 10487 12538
rect 19504 12486 19556 12538
rect 19568 12486 19620 12538
rect 19632 12486 19684 12538
rect 19696 12486 19748 12538
rect 12624 12427 12676 12436
rect 12624 12393 12633 12427
rect 12633 12393 12667 12427
rect 12667 12393 12676 12427
rect 12624 12384 12676 12393
rect 13360 12384 13412 12436
rect 13728 12384 13780 12436
rect 9772 12180 9824 12232
rect 12164 12316 12216 12368
rect 13452 12316 13504 12368
rect 14464 12316 14516 12368
rect 11520 12248 11572 12300
rect 13176 12248 13228 12300
rect 13728 12248 13780 12300
rect 12900 12223 12952 12232
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 12900 12180 12952 12189
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 15568 12180 15620 12232
rect 13268 12112 13320 12164
rect 12440 12044 12492 12096
rect 13452 12044 13504 12096
rect 14556 12044 14608 12096
rect 14648 12044 14700 12096
rect 5612 11942 5664 11994
rect 5676 11942 5728 11994
rect 5740 11942 5792 11994
rect 5804 11942 5856 11994
rect 14874 11942 14926 11994
rect 14938 11942 14990 11994
rect 15002 11942 15054 11994
rect 15066 11942 15118 11994
rect 24135 11942 24187 11994
rect 24199 11942 24251 11994
rect 24263 11942 24315 11994
rect 24327 11942 24379 11994
rect 12900 11840 12952 11892
rect 13268 11883 13320 11892
rect 13268 11849 13277 11883
rect 13277 11849 13311 11883
rect 13311 11849 13320 11883
rect 13268 11840 13320 11849
rect 14096 11840 14148 11892
rect 11060 11772 11112 11824
rect 12716 11704 12768 11756
rect 15108 11704 15160 11756
rect 9680 11568 9732 11620
rect 10876 11636 10928 11688
rect 10968 11636 11020 11688
rect 12256 11679 12308 11688
rect 12256 11645 12265 11679
rect 12265 11645 12299 11679
rect 12299 11645 12308 11679
rect 12256 11636 12308 11645
rect 13084 11636 13136 11688
rect 13360 11636 13412 11688
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 14648 11679 14700 11688
rect 14648 11645 14657 11679
rect 14657 11645 14691 11679
rect 14691 11645 14700 11679
rect 14648 11636 14700 11645
rect 16120 11636 16172 11688
rect 14464 11568 14516 11620
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 10692 11500 10744 11509
rect 14280 11543 14332 11552
rect 14280 11509 14289 11543
rect 14289 11509 14323 11543
rect 14323 11509 14332 11543
rect 14280 11500 14332 11509
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 10243 11398 10295 11450
rect 10307 11398 10359 11450
rect 10371 11398 10423 11450
rect 10435 11398 10487 11450
rect 19504 11398 19556 11450
rect 19568 11398 19620 11450
rect 19632 11398 19684 11450
rect 19696 11398 19748 11450
rect 11520 11339 11572 11348
rect 11520 11305 11529 11339
rect 11529 11305 11563 11339
rect 11563 11305 11572 11339
rect 11520 11296 11572 11305
rect 12716 11339 12768 11348
rect 12716 11305 12725 11339
rect 12725 11305 12759 11339
rect 12759 11305 12768 11339
rect 12716 11296 12768 11305
rect 12992 11296 13044 11348
rect 16120 11339 16172 11348
rect 16120 11305 16129 11339
rect 16129 11305 16163 11339
rect 16163 11305 16172 11339
rect 16120 11296 16172 11305
rect 10692 11228 10744 11280
rect 10968 11228 11020 11280
rect 9772 11160 9824 11212
rect 12440 11228 12492 11280
rect 14648 11228 14700 11280
rect 11980 11160 12032 11212
rect 13820 11203 13872 11212
rect 13544 11092 13596 11144
rect 13820 11169 13829 11203
rect 13829 11169 13863 11203
rect 13863 11169 13872 11203
rect 13820 11160 13872 11169
rect 14556 11160 14608 11212
rect 14648 11092 14700 11144
rect 12348 11024 12400 11076
rect 9680 10999 9732 11008
rect 9680 10965 9689 10999
rect 9689 10965 9723 10999
rect 9723 10965 9732 10999
rect 9680 10956 9732 10965
rect 13360 10999 13412 11008
rect 13360 10965 13369 10999
rect 13369 10965 13403 10999
rect 13403 10965 13412 10999
rect 13360 10956 13412 10965
rect 5612 10854 5664 10906
rect 5676 10854 5728 10906
rect 5740 10854 5792 10906
rect 5804 10854 5856 10906
rect 14874 10854 14926 10906
rect 14938 10854 14990 10906
rect 15002 10854 15054 10906
rect 15066 10854 15118 10906
rect 24135 10854 24187 10906
rect 24199 10854 24251 10906
rect 24263 10854 24315 10906
rect 24327 10854 24379 10906
rect 9956 10795 10008 10804
rect 9956 10761 9965 10795
rect 9965 10761 9999 10795
rect 9999 10761 10008 10795
rect 9956 10752 10008 10761
rect 10968 10795 11020 10804
rect 10968 10761 10977 10795
rect 10977 10761 11011 10795
rect 11011 10761 11020 10795
rect 10968 10752 11020 10761
rect 12256 10752 12308 10804
rect 12532 10795 12584 10804
rect 12532 10761 12541 10795
rect 12541 10761 12575 10795
rect 12575 10761 12584 10795
rect 12532 10752 12584 10761
rect 13360 10752 13412 10804
rect 13820 10752 13872 10804
rect 14280 10795 14332 10804
rect 14280 10761 14289 10795
rect 14289 10761 14323 10795
rect 14323 10761 14332 10795
rect 14280 10752 14332 10761
rect 14648 10752 14700 10804
rect 11060 10684 11112 10736
rect 9680 10548 9732 10600
rect 10600 10480 10652 10532
rect 11520 10548 11572 10600
rect 13544 10616 13596 10668
rect 15384 10684 15436 10736
rect 10968 10455 11020 10464
rect 10968 10421 10998 10455
rect 10998 10421 11020 10455
rect 12164 10455 12216 10464
rect 10968 10412 11020 10421
rect 12164 10421 12173 10455
rect 12173 10421 12207 10455
rect 12207 10421 12216 10455
rect 12164 10412 12216 10421
rect 14188 10548 14240 10600
rect 16120 10616 16172 10668
rect 13820 10480 13872 10532
rect 14372 10480 14424 10532
rect 13912 10412 13964 10464
rect 14096 10455 14148 10464
rect 14096 10421 14105 10455
rect 14105 10421 14139 10455
rect 14139 10421 14148 10455
rect 14096 10412 14148 10421
rect 14188 10412 14240 10464
rect 15568 10480 15620 10532
rect 10243 10310 10295 10362
rect 10307 10310 10359 10362
rect 10371 10310 10423 10362
rect 10435 10310 10487 10362
rect 19504 10310 19556 10362
rect 19568 10310 19620 10362
rect 19632 10310 19684 10362
rect 19696 10310 19748 10362
rect 10600 10208 10652 10260
rect 16120 10251 16172 10260
rect 16120 10217 16129 10251
rect 16129 10217 16163 10251
rect 16163 10217 16172 10251
rect 16120 10208 16172 10217
rect 10968 10140 11020 10192
rect 10140 10072 10192 10124
rect 11980 10072 12032 10124
rect 9772 10004 9824 10056
rect 12164 10072 12216 10124
rect 14188 10072 14240 10124
rect 13820 9979 13872 9988
rect 13820 9945 13829 9979
rect 13829 9945 13863 9979
rect 13863 9945 13872 9979
rect 14648 10004 14700 10056
rect 13820 9936 13872 9945
rect 11428 9911 11480 9920
rect 11428 9877 11437 9911
rect 11437 9877 11471 9911
rect 11471 9877 11480 9911
rect 11428 9868 11480 9877
rect 11888 9911 11940 9920
rect 11888 9877 11897 9911
rect 11897 9877 11931 9911
rect 11931 9877 11940 9911
rect 11888 9868 11940 9877
rect 5612 9766 5664 9818
rect 5676 9766 5728 9818
rect 5740 9766 5792 9818
rect 5804 9766 5856 9818
rect 14874 9766 14926 9818
rect 14938 9766 14990 9818
rect 15002 9766 15054 9818
rect 15066 9766 15118 9818
rect 24135 9766 24187 9818
rect 24199 9766 24251 9818
rect 24263 9766 24315 9818
rect 24327 9766 24379 9818
rect 12164 9707 12216 9716
rect 12164 9673 12173 9707
rect 12173 9673 12207 9707
rect 12207 9673 12216 9707
rect 12164 9664 12216 9673
rect 14280 9664 14332 9716
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 11520 9528 11572 9580
rect 13912 9528 13964 9580
rect 15292 9571 15344 9580
rect 15292 9537 15301 9571
rect 15301 9537 15335 9571
rect 15335 9537 15344 9571
rect 15292 9528 15344 9537
rect 12256 9503 12308 9512
rect 12256 9469 12265 9503
rect 12265 9469 12299 9503
rect 12299 9469 12308 9503
rect 12256 9460 12308 9469
rect 13820 9503 13872 9512
rect 10876 9392 10928 9444
rect 12072 9392 12124 9444
rect 13820 9469 13829 9503
rect 13829 9469 13863 9503
rect 13863 9469 13872 9503
rect 13820 9460 13872 9469
rect 14464 9392 14516 9444
rect 15200 9460 15252 9512
rect 16212 9392 16264 9444
rect 16120 9367 16172 9376
rect 16120 9333 16129 9367
rect 16129 9333 16163 9367
rect 16163 9333 16172 9367
rect 16120 9324 16172 9333
rect 10243 9222 10295 9274
rect 10307 9222 10359 9274
rect 10371 9222 10423 9274
rect 10435 9222 10487 9274
rect 19504 9222 19556 9274
rect 19568 9222 19620 9274
rect 19632 9222 19684 9274
rect 19696 9222 19748 9274
rect 10140 9120 10192 9172
rect 10968 9163 11020 9172
rect 10968 9129 10977 9163
rect 10977 9129 11011 9163
rect 11011 9129 11020 9163
rect 10968 9120 11020 9129
rect 11520 9120 11572 9172
rect 16120 9052 16172 9104
rect 10600 8984 10652 9036
rect 11428 8984 11480 9036
rect 11796 8984 11848 9036
rect 14648 8984 14700 9036
rect 10140 8848 10192 8900
rect 13728 8848 13780 8900
rect 11520 8823 11572 8832
rect 11520 8789 11529 8823
rect 11529 8789 11563 8823
rect 11563 8789 11572 8823
rect 11520 8780 11572 8789
rect 16120 8823 16172 8832
rect 16120 8789 16129 8823
rect 16129 8789 16163 8823
rect 16163 8789 16172 8823
rect 16120 8780 16172 8789
rect 5612 8678 5664 8730
rect 5676 8678 5728 8730
rect 5740 8678 5792 8730
rect 5804 8678 5856 8730
rect 14874 8678 14926 8730
rect 14938 8678 14990 8730
rect 15002 8678 15054 8730
rect 15066 8678 15118 8730
rect 24135 8678 24187 8730
rect 24199 8678 24251 8730
rect 24263 8678 24315 8730
rect 24327 8678 24379 8730
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 11520 8576 11572 8628
rect 15292 8483 15344 8492
rect 11888 8372 11940 8424
rect 12072 8415 12124 8424
rect 12072 8381 12081 8415
rect 12081 8381 12115 8415
rect 12115 8381 12124 8415
rect 12072 8372 12124 8381
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 15292 8449 15301 8483
rect 15301 8449 15335 8483
rect 15335 8449 15344 8483
rect 15292 8440 15344 8449
rect 12256 8372 12308 8381
rect 14556 8415 14608 8424
rect 14556 8381 14565 8415
rect 14565 8381 14599 8415
rect 14599 8381 14608 8415
rect 14556 8372 14608 8381
rect 15200 8415 15252 8424
rect 15200 8381 15209 8415
rect 15209 8381 15243 8415
rect 15243 8381 15252 8415
rect 15200 8372 15252 8381
rect 16120 8372 16172 8424
rect 10243 8134 10295 8186
rect 10307 8134 10359 8186
rect 10371 8134 10423 8186
rect 10435 8134 10487 8186
rect 19504 8134 19556 8186
rect 19568 8134 19620 8186
rect 19632 8134 19684 8186
rect 19696 8134 19748 8186
rect 12348 8032 12400 8084
rect 12164 7964 12216 8016
rect 14740 7964 14792 8016
rect 12532 7939 12584 7948
rect 9772 7828 9824 7880
rect 10600 7871 10652 7880
rect 10600 7837 10609 7871
rect 10609 7837 10643 7871
rect 10643 7837 10652 7871
rect 10600 7828 10652 7837
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 12532 7905 12541 7939
rect 12541 7905 12575 7939
rect 12575 7905 12584 7939
rect 12532 7896 12584 7905
rect 12808 7939 12860 7948
rect 12808 7905 12817 7939
rect 12817 7905 12851 7939
rect 12851 7905 12860 7939
rect 12808 7896 12860 7905
rect 13820 7828 13872 7880
rect 12256 7760 12308 7812
rect 13452 7760 13504 7812
rect 10876 7692 10928 7744
rect 12072 7735 12124 7744
rect 12072 7701 12081 7735
rect 12081 7701 12115 7735
rect 12115 7701 12124 7735
rect 12072 7692 12124 7701
rect 12348 7692 12400 7744
rect 15384 7692 15436 7744
rect 5612 7590 5664 7642
rect 5676 7590 5728 7642
rect 5740 7590 5792 7642
rect 5804 7590 5856 7642
rect 14874 7590 14926 7642
rect 14938 7590 14990 7642
rect 15002 7590 15054 7642
rect 15066 7590 15118 7642
rect 24135 7590 24187 7642
rect 24199 7590 24251 7642
rect 24263 7590 24315 7642
rect 24327 7590 24379 7642
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 12256 7531 12308 7540
rect 12256 7497 12265 7531
rect 12265 7497 12299 7531
rect 12299 7497 12308 7531
rect 12256 7488 12308 7497
rect 14740 7531 14792 7540
rect 14740 7497 14749 7531
rect 14749 7497 14783 7531
rect 14783 7497 14792 7531
rect 14740 7488 14792 7497
rect 10876 7327 10928 7336
rect 10876 7293 10894 7327
rect 10894 7293 10928 7327
rect 10876 7284 10928 7293
rect 11060 7284 11112 7336
rect 13820 7352 13872 7404
rect 13912 7352 13964 7404
rect 15108 7420 15160 7472
rect 13452 7284 13504 7336
rect 10600 7216 10652 7268
rect 12900 7216 12952 7268
rect 13360 7216 13412 7268
rect 15108 7284 15160 7336
rect 15384 7327 15436 7336
rect 15384 7293 15393 7327
rect 15393 7293 15427 7327
rect 15427 7293 15436 7327
rect 15384 7284 15436 7293
rect 14556 7216 14608 7268
rect 12716 7148 12768 7200
rect 14464 7148 14516 7200
rect 15016 7148 15068 7200
rect 10243 7046 10295 7098
rect 10307 7046 10359 7098
rect 10371 7046 10423 7098
rect 10435 7046 10487 7098
rect 19504 7046 19556 7098
rect 19568 7046 19620 7098
rect 19632 7046 19684 7098
rect 19696 7046 19748 7098
rect 12072 6876 12124 6928
rect 10692 6808 10744 6860
rect 10968 6808 11020 6860
rect 12164 6808 12216 6860
rect 12440 6851 12492 6860
rect 12440 6817 12449 6851
rect 12449 6817 12483 6851
rect 12483 6817 12492 6851
rect 12440 6808 12492 6817
rect 12348 6740 12400 6792
rect 12716 6740 12768 6792
rect 11888 6672 11940 6724
rect 13268 6808 13320 6860
rect 13544 6808 13596 6860
rect 13636 6672 13688 6724
rect 11060 6604 11112 6656
rect 11704 6604 11756 6656
rect 12532 6604 12584 6656
rect 13360 6604 13412 6656
rect 15016 6808 15068 6860
rect 14740 6740 14792 6792
rect 14464 6604 14516 6656
rect 15384 6647 15436 6656
rect 15384 6613 15393 6647
rect 15393 6613 15427 6647
rect 15427 6613 15436 6647
rect 15384 6604 15436 6613
rect 5612 6502 5664 6554
rect 5676 6502 5728 6554
rect 5740 6502 5792 6554
rect 5804 6502 5856 6554
rect 14874 6502 14926 6554
rect 14938 6502 14990 6554
rect 15002 6502 15054 6554
rect 15066 6502 15118 6554
rect 24135 6502 24187 6554
rect 24199 6502 24251 6554
rect 24263 6502 24315 6554
rect 24327 6502 24379 6554
rect 11888 6400 11940 6452
rect 12440 6400 12492 6452
rect 13452 6400 13504 6452
rect 10140 6239 10192 6248
rect 10140 6205 10149 6239
rect 10149 6205 10183 6239
rect 10183 6205 10192 6239
rect 10140 6196 10192 6205
rect 11520 6196 11572 6248
rect 12072 6196 12124 6248
rect 12716 6239 12768 6248
rect 12716 6205 12725 6239
rect 12725 6205 12759 6239
rect 12759 6205 12768 6239
rect 13360 6239 13412 6248
rect 12716 6196 12768 6205
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 13820 6239 13872 6248
rect 13820 6205 13829 6239
rect 13829 6205 13863 6239
rect 13863 6205 13872 6239
rect 13820 6196 13872 6205
rect 15384 6196 15436 6248
rect 11060 6128 11112 6180
rect 12348 6171 12400 6180
rect 12348 6137 12357 6171
rect 12357 6137 12391 6171
rect 12391 6137 12400 6171
rect 12348 6128 12400 6137
rect 10692 6060 10744 6112
rect 12256 6060 12308 6112
rect 13268 6128 13320 6180
rect 16396 6128 16448 6180
rect 14924 6060 14976 6112
rect 10243 5958 10295 6010
rect 10307 5958 10359 6010
rect 10371 5958 10423 6010
rect 10435 5958 10487 6010
rect 19504 5958 19556 6010
rect 19568 5958 19620 6010
rect 19632 5958 19684 6010
rect 19696 5958 19748 6010
rect 12164 5856 12216 5908
rect 13820 5856 13872 5908
rect 14740 5856 14792 5908
rect 10600 5788 10652 5840
rect 11520 5831 11572 5840
rect 11520 5797 11529 5831
rect 11529 5797 11563 5831
rect 11563 5797 11572 5831
rect 11520 5788 11572 5797
rect 12348 5788 12400 5840
rect 10048 5652 10100 5704
rect 11152 5720 11204 5772
rect 11980 5720 12032 5772
rect 13360 5788 13412 5840
rect 12900 5720 12952 5772
rect 12992 5720 13044 5772
rect 13912 5720 13964 5772
rect 14924 5763 14976 5772
rect 14924 5729 14933 5763
rect 14933 5729 14967 5763
rect 14967 5729 14976 5763
rect 14924 5720 14976 5729
rect 14464 5584 14516 5636
rect 13544 5516 13596 5568
rect 15660 5516 15712 5568
rect 5612 5414 5664 5466
rect 5676 5414 5728 5466
rect 5740 5414 5792 5466
rect 5804 5414 5856 5466
rect 14874 5414 14926 5466
rect 14938 5414 14990 5466
rect 15002 5414 15054 5466
rect 15066 5414 15118 5466
rect 24135 5414 24187 5466
rect 24199 5414 24251 5466
rect 24263 5414 24315 5466
rect 24327 5414 24379 5466
rect 12348 5312 12400 5364
rect 12808 5312 12860 5364
rect 12256 5176 12308 5228
rect 12532 5219 12584 5228
rect 12532 5185 12541 5219
rect 12541 5185 12575 5219
rect 12575 5185 12584 5219
rect 12532 5176 12584 5185
rect 11520 5108 11572 5160
rect 12348 5108 12400 5160
rect 12624 5151 12676 5160
rect 12624 5117 12633 5151
rect 12633 5117 12667 5151
rect 12667 5117 12676 5151
rect 12624 5108 12676 5117
rect 12716 5151 12768 5160
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 12716 5108 12768 5117
rect 13636 5108 13688 5160
rect 14004 5176 14056 5228
rect 13820 5151 13872 5160
rect 13820 5117 13829 5151
rect 13829 5117 13863 5151
rect 13863 5117 13872 5151
rect 13820 5108 13872 5117
rect 14464 5151 14516 5160
rect 14464 5117 14473 5151
rect 14473 5117 14507 5151
rect 14507 5117 14516 5151
rect 14464 5108 14516 5117
rect 15936 5151 15988 5160
rect 15936 5117 15945 5151
rect 15945 5117 15979 5151
rect 15979 5117 15988 5151
rect 15936 5108 15988 5117
rect 11060 5015 11112 5024
rect 11060 4981 11069 5015
rect 11069 4981 11103 5015
rect 11103 4981 11112 5015
rect 11060 4972 11112 4981
rect 13544 4972 13596 5024
rect 16212 4972 16264 5024
rect 10243 4870 10295 4922
rect 10307 4870 10359 4922
rect 10371 4870 10423 4922
rect 10435 4870 10487 4922
rect 19504 4870 19556 4922
rect 19568 4870 19620 4922
rect 19632 4870 19684 4922
rect 19696 4870 19748 4922
rect 12716 4811 12768 4820
rect 12716 4777 12718 4811
rect 12718 4777 12752 4811
rect 12752 4777 12768 4811
rect 11060 4700 11112 4752
rect 12716 4768 12768 4777
rect 12900 4768 12952 4820
rect 13912 4768 13964 4820
rect 16212 4811 16264 4820
rect 16212 4777 16221 4811
rect 16221 4777 16255 4811
rect 16255 4777 16264 4811
rect 16212 4768 16264 4777
rect 12164 4700 12216 4752
rect 12348 4700 12400 4752
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 10600 4632 10652 4684
rect 12532 4675 12584 4684
rect 12532 4641 12541 4675
rect 12541 4641 12575 4675
rect 12575 4641 12584 4675
rect 12532 4632 12584 4641
rect 12624 4675 12676 4684
rect 12624 4641 12633 4675
rect 12633 4641 12667 4675
rect 12667 4641 12676 4675
rect 12624 4632 12676 4641
rect 12348 4564 12400 4616
rect 14004 4632 14056 4684
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 17868 4632 17920 4684
rect 14372 4564 14424 4616
rect 16396 4607 16448 4616
rect 16396 4573 16405 4607
rect 16405 4573 16439 4607
rect 16439 4573 16448 4607
rect 16396 4564 16448 4573
rect 13268 4539 13320 4548
rect 13268 4505 13277 4539
rect 13277 4505 13311 4539
rect 13311 4505 13320 4539
rect 13268 4496 13320 4505
rect 9956 4471 10008 4480
rect 9956 4437 9965 4471
rect 9965 4437 9999 4471
rect 9999 4437 10008 4471
rect 9956 4428 10008 4437
rect 15292 4428 15344 4480
rect 15844 4471 15896 4480
rect 15844 4437 15853 4471
rect 15853 4437 15887 4471
rect 15887 4437 15896 4471
rect 15844 4428 15896 4437
rect 5612 4326 5664 4378
rect 5676 4326 5728 4378
rect 5740 4326 5792 4378
rect 5804 4326 5856 4378
rect 14874 4326 14926 4378
rect 14938 4326 14990 4378
rect 15002 4326 15054 4378
rect 15066 4326 15118 4378
rect 24135 4326 24187 4378
rect 24199 4326 24251 4378
rect 24263 4326 24315 4378
rect 24327 4326 24379 4378
rect 12532 4224 12584 4276
rect 14372 4267 14424 4276
rect 14372 4233 14381 4267
rect 14381 4233 14415 4267
rect 14415 4233 14424 4267
rect 14372 4224 14424 4233
rect 15936 4224 15988 4276
rect 11152 4063 11204 4072
rect 11152 4029 11161 4063
rect 11161 4029 11195 4063
rect 11195 4029 11204 4063
rect 11152 4020 11204 4029
rect 12164 4063 12216 4072
rect 12164 4029 12173 4063
rect 12173 4029 12207 4063
rect 12207 4029 12216 4063
rect 12164 4020 12216 4029
rect 10600 3952 10652 4004
rect 11796 3952 11848 4004
rect 12808 4156 12860 4208
rect 12624 4088 12676 4140
rect 12900 4020 12952 4072
rect 13820 4020 13872 4072
rect 15292 4063 15344 4072
rect 15292 4029 15326 4063
rect 15326 4029 15344 4063
rect 15292 4020 15344 4029
rect 12808 3952 12860 4004
rect 13728 3952 13780 4004
rect 12348 3884 12400 3936
rect 12992 3884 13044 3936
rect 10243 3782 10295 3834
rect 10307 3782 10359 3834
rect 10371 3782 10423 3834
rect 10435 3782 10487 3834
rect 19504 3782 19556 3834
rect 19568 3782 19620 3834
rect 19632 3782 19684 3834
rect 19696 3782 19748 3834
rect 13268 3680 13320 3732
rect 14740 3680 14792 3732
rect 15844 3680 15896 3732
rect 9956 3612 10008 3664
rect 10692 3544 10744 3596
rect 13544 3587 13596 3596
rect 13544 3553 13562 3587
rect 13562 3553 13596 3587
rect 13820 3587 13872 3596
rect 13544 3544 13596 3553
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 13820 3544 13872 3553
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 27896 3476 27948 3528
rect 12900 3340 12952 3392
rect 5612 3238 5664 3290
rect 5676 3238 5728 3290
rect 5740 3238 5792 3290
rect 5804 3238 5856 3290
rect 14874 3238 14926 3290
rect 14938 3238 14990 3290
rect 15002 3238 15054 3290
rect 15066 3238 15118 3290
rect 24135 3238 24187 3290
rect 24199 3238 24251 3290
rect 24263 3238 24315 3290
rect 24327 3238 24379 3290
rect 12256 3136 12308 3188
rect 17868 3136 17920 3188
rect 27896 3179 27948 3188
rect 27896 3145 27905 3179
rect 27905 3145 27939 3179
rect 27939 3145 27948 3179
rect 27896 3136 27948 3145
rect 12624 3000 12676 3052
rect 12532 2932 12584 2984
rect 13268 2932 13320 2984
rect 14372 2932 14424 2984
rect 20720 2932 20772 2984
rect 27344 2932 27396 2984
rect 10243 2694 10295 2746
rect 10307 2694 10359 2746
rect 10371 2694 10423 2746
rect 10435 2694 10487 2746
rect 19504 2694 19556 2746
rect 19568 2694 19620 2746
rect 19632 2694 19684 2746
rect 19696 2694 19748 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 20720 2635 20772 2644
rect 20720 2601 20729 2635
rect 20729 2601 20763 2635
rect 20763 2601 20772 2635
rect 20720 2592 20772 2601
rect 27344 2635 27396 2644
rect 27344 2601 27353 2635
rect 27353 2601 27387 2635
rect 27387 2601 27396 2635
rect 27344 2592 27396 2601
rect 480 2456 532 2508
rect 20720 2456 20772 2508
rect 27160 2499 27212 2508
rect 27160 2465 27169 2499
rect 27169 2465 27203 2499
rect 27203 2465 27212 2499
rect 27160 2456 27212 2465
rect 5612 2150 5664 2202
rect 5676 2150 5728 2202
rect 5740 2150 5792 2202
rect 5804 2150 5856 2202
rect 14874 2150 14926 2202
rect 14938 2150 14990 2202
rect 15002 2150 15054 2202
rect 15066 2150 15118 2202
rect 24135 2150 24187 2202
rect 24199 2150 24251 2202
rect 24263 2150 24315 2202
rect 24327 2150 24379 2202
<< metal2 >>
rect 9218 31368 9274 32168
rect 19338 31368 19394 32168
rect 29458 31368 29514 32168
rect 1398 30016 1454 30025
rect 1398 29951 1454 29960
rect 1412 29714 1440 29951
rect 9232 29714 9260 31368
rect 10217 29948 10513 29968
rect 10273 29946 10297 29948
rect 10353 29946 10377 29948
rect 10433 29946 10457 29948
rect 10295 29894 10297 29946
rect 10359 29894 10371 29946
rect 10433 29894 10435 29946
rect 10273 29892 10297 29894
rect 10353 29892 10377 29894
rect 10433 29892 10457 29894
rect 10217 29872 10513 29892
rect 19352 29714 19380 31368
rect 19478 29948 19774 29968
rect 19534 29946 19558 29948
rect 19614 29946 19638 29948
rect 19694 29946 19718 29948
rect 19556 29894 19558 29946
rect 19620 29894 19632 29946
rect 19694 29894 19696 29946
rect 19534 29892 19558 29894
rect 19614 29892 19638 29894
rect 19694 29892 19718 29894
rect 19478 29872 19774 29892
rect 29472 29782 29500 31368
rect 29460 29776 29512 29782
rect 29460 29718 29512 29724
rect 1400 29708 1452 29714
rect 1400 29650 1452 29656
rect 9220 29708 9272 29714
rect 9220 29650 9272 29656
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 1584 29504 1636 29510
rect 1584 29446 1636 29452
rect 9772 29504 9824 29510
rect 9772 29446 9824 29452
rect 14740 29504 14792 29510
rect 14740 29446 14792 29452
rect 1398 15056 1454 15065
rect 1596 15026 1624 29446
rect 5586 29404 5882 29424
rect 5642 29402 5666 29404
rect 5722 29402 5746 29404
rect 5802 29402 5826 29404
rect 5664 29350 5666 29402
rect 5728 29350 5740 29402
rect 5802 29350 5804 29402
rect 5642 29348 5666 29350
rect 5722 29348 5746 29350
rect 5802 29348 5826 29350
rect 5586 29328 5882 29348
rect 5586 28316 5882 28336
rect 5642 28314 5666 28316
rect 5722 28314 5746 28316
rect 5802 28314 5826 28316
rect 5664 28262 5666 28314
rect 5728 28262 5740 28314
rect 5802 28262 5804 28314
rect 5642 28260 5666 28262
rect 5722 28260 5746 28262
rect 5802 28260 5826 28262
rect 5586 28240 5882 28260
rect 5586 27228 5882 27248
rect 5642 27226 5666 27228
rect 5722 27226 5746 27228
rect 5802 27226 5826 27228
rect 5664 27174 5666 27226
rect 5728 27174 5740 27226
rect 5802 27174 5804 27226
rect 5642 27172 5666 27174
rect 5722 27172 5746 27174
rect 5802 27172 5826 27174
rect 5586 27152 5882 27172
rect 5586 26140 5882 26160
rect 5642 26138 5666 26140
rect 5722 26138 5746 26140
rect 5802 26138 5826 26140
rect 5664 26086 5666 26138
rect 5728 26086 5740 26138
rect 5802 26086 5804 26138
rect 5642 26084 5666 26086
rect 5722 26084 5746 26086
rect 5802 26084 5826 26086
rect 5586 26064 5882 26084
rect 5586 25052 5882 25072
rect 5642 25050 5666 25052
rect 5722 25050 5746 25052
rect 5802 25050 5826 25052
rect 5664 24998 5666 25050
rect 5728 24998 5740 25050
rect 5802 24998 5804 25050
rect 5642 24996 5666 24998
rect 5722 24996 5746 24998
rect 5802 24996 5826 24998
rect 5586 24976 5882 24996
rect 5586 23964 5882 23984
rect 5642 23962 5666 23964
rect 5722 23962 5746 23964
rect 5802 23962 5826 23964
rect 5664 23910 5666 23962
rect 5728 23910 5740 23962
rect 5802 23910 5804 23962
rect 5642 23908 5666 23910
rect 5722 23908 5746 23910
rect 5802 23908 5826 23910
rect 5586 23888 5882 23908
rect 5586 22876 5882 22896
rect 5642 22874 5666 22876
rect 5722 22874 5746 22876
rect 5802 22874 5826 22876
rect 5664 22822 5666 22874
rect 5728 22822 5740 22874
rect 5802 22822 5804 22874
rect 5642 22820 5666 22822
rect 5722 22820 5746 22822
rect 5802 22820 5826 22822
rect 5586 22800 5882 22820
rect 5586 21788 5882 21808
rect 5642 21786 5666 21788
rect 5722 21786 5746 21788
rect 5802 21786 5826 21788
rect 5664 21734 5666 21786
rect 5728 21734 5740 21786
rect 5802 21734 5804 21786
rect 5642 21732 5666 21734
rect 5722 21732 5746 21734
rect 5802 21732 5826 21734
rect 5586 21712 5882 21732
rect 5586 20700 5882 20720
rect 5642 20698 5666 20700
rect 5722 20698 5746 20700
rect 5802 20698 5826 20700
rect 5664 20646 5666 20698
rect 5728 20646 5740 20698
rect 5802 20646 5804 20698
rect 5642 20644 5666 20646
rect 5722 20644 5746 20646
rect 5802 20644 5826 20646
rect 5586 20624 5882 20644
rect 5586 19612 5882 19632
rect 5642 19610 5666 19612
rect 5722 19610 5746 19612
rect 5802 19610 5826 19612
rect 5664 19558 5666 19610
rect 5728 19558 5740 19610
rect 5802 19558 5804 19610
rect 5642 19556 5666 19558
rect 5722 19556 5746 19558
rect 5802 19556 5826 19558
rect 5586 19536 5882 19556
rect 5586 18524 5882 18544
rect 5642 18522 5666 18524
rect 5722 18522 5746 18524
rect 5802 18522 5826 18524
rect 5664 18470 5666 18522
rect 5728 18470 5740 18522
rect 5802 18470 5804 18522
rect 5642 18468 5666 18470
rect 5722 18468 5746 18470
rect 5802 18468 5826 18470
rect 5586 18448 5882 18468
rect 5586 17436 5882 17456
rect 5642 17434 5666 17436
rect 5722 17434 5746 17436
rect 5802 17434 5826 17436
rect 5664 17382 5666 17434
rect 5728 17382 5740 17434
rect 5802 17382 5804 17434
rect 5642 17380 5666 17382
rect 5722 17380 5746 17382
rect 5802 17380 5826 17382
rect 5586 17360 5882 17380
rect 5586 16348 5882 16368
rect 5642 16346 5666 16348
rect 5722 16346 5746 16348
rect 5802 16346 5826 16348
rect 5664 16294 5666 16346
rect 5728 16294 5740 16346
rect 5802 16294 5804 16346
rect 5642 16292 5666 16294
rect 5722 16292 5746 16294
rect 5802 16292 5826 16294
rect 5586 16272 5882 16292
rect 5586 15260 5882 15280
rect 5642 15258 5666 15260
rect 5722 15258 5746 15260
rect 5802 15258 5826 15260
rect 5664 15206 5666 15258
rect 5728 15206 5740 15258
rect 5802 15206 5804 15258
rect 5642 15204 5666 15206
rect 5722 15204 5746 15206
rect 5802 15204 5826 15206
rect 5586 15184 5882 15204
rect 1398 14991 1454 15000
rect 1584 15020 1636 15026
rect 1412 14958 1440 14991
rect 1584 14962 1636 14968
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8496 14550 8524 14758
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 5586 14172 5882 14192
rect 5642 14170 5666 14172
rect 5722 14170 5746 14172
rect 5802 14170 5826 14172
rect 5664 14118 5666 14170
rect 5728 14118 5740 14170
rect 5802 14118 5804 14170
rect 5642 14116 5666 14118
rect 5722 14116 5746 14118
rect 5802 14116 5826 14118
rect 5586 14096 5882 14116
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 1596 2650 1624 13330
rect 9784 13326 9812 29446
rect 10217 28860 10513 28880
rect 10273 28858 10297 28860
rect 10353 28858 10377 28860
rect 10433 28858 10457 28860
rect 10295 28806 10297 28858
rect 10359 28806 10371 28858
rect 10433 28806 10435 28858
rect 10273 28804 10297 28806
rect 10353 28804 10377 28806
rect 10433 28804 10457 28806
rect 10217 28784 10513 28804
rect 10217 27772 10513 27792
rect 10273 27770 10297 27772
rect 10353 27770 10377 27772
rect 10433 27770 10457 27772
rect 10295 27718 10297 27770
rect 10359 27718 10371 27770
rect 10433 27718 10435 27770
rect 10273 27716 10297 27718
rect 10353 27716 10377 27718
rect 10433 27716 10457 27718
rect 10217 27696 10513 27716
rect 10217 26684 10513 26704
rect 10273 26682 10297 26684
rect 10353 26682 10377 26684
rect 10433 26682 10457 26684
rect 10295 26630 10297 26682
rect 10359 26630 10371 26682
rect 10433 26630 10435 26682
rect 10273 26628 10297 26630
rect 10353 26628 10377 26630
rect 10433 26628 10457 26630
rect 10217 26608 10513 26628
rect 10217 25596 10513 25616
rect 10273 25594 10297 25596
rect 10353 25594 10377 25596
rect 10433 25594 10457 25596
rect 10295 25542 10297 25594
rect 10359 25542 10371 25594
rect 10433 25542 10435 25594
rect 10273 25540 10297 25542
rect 10353 25540 10377 25542
rect 10433 25540 10457 25542
rect 10217 25520 10513 25540
rect 10217 24508 10513 24528
rect 10273 24506 10297 24508
rect 10353 24506 10377 24508
rect 10433 24506 10457 24508
rect 10295 24454 10297 24506
rect 10359 24454 10371 24506
rect 10433 24454 10435 24506
rect 10273 24452 10297 24454
rect 10353 24452 10377 24454
rect 10433 24452 10457 24454
rect 10217 24432 10513 24452
rect 10217 23420 10513 23440
rect 10273 23418 10297 23420
rect 10353 23418 10377 23420
rect 10433 23418 10457 23420
rect 10295 23366 10297 23418
rect 10359 23366 10371 23418
rect 10433 23366 10435 23418
rect 10273 23364 10297 23366
rect 10353 23364 10377 23366
rect 10433 23364 10457 23366
rect 10217 23344 10513 23364
rect 10217 22332 10513 22352
rect 10273 22330 10297 22332
rect 10353 22330 10377 22332
rect 10433 22330 10457 22332
rect 10295 22278 10297 22330
rect 10359 22278 10371 22330
rect 10433 22278 10435 22330
rect 10273 22276 10297 22278
rect 10353 22276 10377 22278
rect 10433 22276 10457 22278
rect 10217 22256 10513 22276
rect 10217 21244 10513 21264
rect 10273 21242 10297 21244
rect 10353 21242 10377 21244
rect 10433 21242 10457 21244
rect 10295 21190 10297 21242
rect 10359 21190 10371 21242
rect 10433 21190 10435 21242
rect 10273 21188 10297 21190
rect 10353 21188 10377 21190
rect 10433 21188 10457 21190
rect 10217 21168 10513 21188
rect 10217 20156 10513 20176
rect 10273 20154 10297 20156
rect 10353 20154 10377 20156
rect 10433 20154 10457 20156
rect 10295 20102 10297 20154
rect 10359 20102 10371 20154
rect 10433 20102 10435 20154
rect 10273 20100 10297 20102
rect 10353 20100 10377 20102
rect 10433 20100 10457 20102
rect 10217 20080 10513 20100
rect 10217 19068 10513 19088
rect 10273 19066 10297 19068
rect 10353 19066 10377 19068
rect 10433 19066 10457 19068
rect 10295 19014 10297 19066
rect 10359 19014 10371 19066
rect 10433 19014 10435 19066
rect 10273 19012 10297 19014
rect 10353 19012 10377 19014
rect 10433 19012 10457 19014
rect 10217 18992 10513 19012
rect 10217 17980 10513 18000
rect 10273 17978 10297 17980
rect 10353 17978 10377 17980
rect 10433 17978 10457 17980
rect 10295 17926 10297 17978
rect 10359 17926 10371 17978
rect 10433 17926 10435 17978
rect 10273 17924 10297 17926
rect 10353 17924 10377 17926
rect 10433 17924 10457 17926
rect 10217 17904 10513 17924
rect 10217 16892 10513 16912
rect 10273 16890 10297 16892
rect 10353 16890 10377 16892
rect 10433 16890 10457 16892
rect 10295 16838 10297 16890
rect 10359 16838 10371 16890
rect 10433 16838 10435 16890
rect 10273 16836 10297 16838
rect 10353 16836 10377 16838
rect 10433 16836 10457 16838
rect 10217 16816 10513 16836
rect 10217 15804 10513 15824
rect 10273 15802 10297 15804
rect 10353 15802 10377 15804
rect 10433 15802 10457 15804
rect 10295 15750 10297 15802
rect 10359 15750 10371 15802
rect 10433 15750 10435 15802
rect 10273 15748 10297 15750
rect 10353 15748 10377 15750
rect 10433 15748 10457 15750
rect 10217 15728 10513 15748
rect 14752 15570 14780 29446
rect 14848 29404 15144 29424
rect 14904 29402 14928 29404
rect 14984 29402 15008 29404
rect 15064 29402 15088 29404
rect 14926 29350 14928 29402
rect 14990 29350 15002 29402
rect 15064 29350 15066 29402
rect 14904 29348 14928 29350
rect 14984 29348 15008 29350
rect 15064 29348 15088 29350
rect 14848 29328 15144 29348
rect 24109 29404 24405 29424
rect 24165 29402 24189 29404
rect 24245 29402 24269 29404
rect 24325 29402 24349 29404
rect 24187 29350 24189 29402
rect 24251 29350 24263 29402
rect 24325 29350 24327 29402
rect 24165 29348 24189 29350
rect 24245 29348 24269 29350
rect 24325 29348 24349 29350
rect 24109 29328 24405 29348
rect 19478 28860 19774 28880
rect 19534 28858 19558 28860
rect 19614 28858 19638 28860
rect 19694 28858 19718 28860
rect 19556 28806 19558 28858
rect 19620 28806 19632 28858
rect 19694 28806 19696 28858
rect 19534 28804 19558 28806
rect 19614 28804 19638 28806
rect 19694 28804 19718 28806
rect 19478 28784 19774 28804
rect 14848 28316 15144 28336
rect 14904 28314 14928 28316
rect 14984 28314 15008 28316
rect 15064 28314 15088 28316
rect 14926 28262 14928 28314
rect 14990 28262 15002 28314
rect 15064 28262 15066 28314
rect 14904 28260 14928 28262
rect 14984 28260 15008 28262
rect 15064 28260 15088 28262
rect 14848 28240 15144 28260
rect 24109 28316 24405 28336
rect 24165 28314 24189 28316
rect 24245 28314 24269 28316
rect 24325 28314 24349 28316
rect 24187 28262 24189 28314
rect 24251 28262 24263 28314
rect 24325 28262 24327 28314
rect 24165 28260 24189 28262
rect 24245 28260 24269 28262
rect 24325 28260 24349 28262
rect 24109 28240 24405 28260
rect 19478 27772 19774 27792
rect 19534 27770 19558 27772
rect 19614 27770 19638 27772
rect 19694 27770 19718 27772
rect 19556 27718 19558 27770
rect 19620 27718 19632 27770
rect 19694 27718 19696 27770
rect 19534 27716 19558 27718
rect 19614 27716 19638 27718
rect 19694 27716 19718 27718
rect 19478 27696 19774 27716
rect 14848 27228 15144 27248
rect 14904 27226 14928 27228
rect 14984 27226 15008 27228
rect 15064 27226 15088 27228
rect 14926 27174 14928 27226
rect 14990 27174 15002 27226
rect 15064 27174 15066 27226
rect 14904 27172 14928 27174
rect 14984 27172 15008 27174
rect 15064 27172 15088 27174
rect 14848 27152 15144 27172
rect 24109 27228 24405 27248
rect 24165 27226 24189 27228
rect 24245 27226 24269 27228
rect 24325 27226 24349 27228
rect 24187 27174 24189 27226
rect 24251 27174 24263 27226
rect 24325 27174 24327 27226
rect 24165 27172 24189 27174
rect 24245 27172 24269 27174
rect 24325 27172 24349 27174
rect 24109 27152 24405 27172
rect 19478 26684 19774 26704
rect 19534 26682 19558 26684
rect 19614 26682 19638 26684
rect 19694 26682 19718 26684
rect 19556 26630 19558 26682
rect 19620 26630 19632 26682
rect 19694 26630 19696 26682
rect 19534 26628 19558 26630
rect 19614 26628 19638 26630
rect 19694 26628 19718 26630
rect 19478 26608 19774 26628
rect 14848 26140 15144 26160
rect 14904 26138 14928 26140
rect 14984 26138 15008 26140
rect 15064 26138 15088 26140
rect 14926 26086 14928 26138
rect 14990 26086 15002 26138
rect 15064 26086 15066 26138
rect 14904 26084 14928 26086
rect 14984 26084 15008 26086
rect 15064 26084 15088 26086
rect 14848 26064 15144 26084
rect 24109 26140 24405 26160
rect 24165 26138 24189 26140
rect 24245 26138 24269 26140
rect 24325 26138 24349 26140
rect 24187 26086 24189 26138
rect 24251 26086 24263 26138
rect 24325 26086 24327 26138
rect 24165 26084 24189 26086
rect 24245 26084 24269 26086
rect 24325 26084 24349 26086
rect 24109 26064 24405 26084
rect 19478 25596 19774 25616
rect 19534 25594 19558 25596
rect 19614 25594 19638 25596
rect 19694 25594 19718 25596
rect 19556 25542 19558 25594
rect 19620 25542 19632 25594
rect 19694 25542 19696 25594
rect 19534 25540 19558 25542
rect 19614 25540 19638 25542
rect 19694 25540 19718 25542
rect 19478 25520 19774 25540
rect 14848 25052 15144 25072
rect 14904 25050 14928 25052
rect 14984 25050 15008 25052
rect 15064 25050 15088 25052
rect 14926 24998 14928 25050
rect 14990 24998 15002 25050
rect 15064 24998 15066 25050
rect 14904 24996 14928 24998
rect 14984 24996 15008 24998
rect 15064 24996 15088 24998
rect 14848 24976 15144 24996
rect 24109 25052 24405 25072
rect 24165 25050 24189 25052
rect 24245 25050 24269 25052
rect 24325 25050 24349 25052
rect 24187 24998 24189 25050
rect 24251 24998 24263 25050
rect 24325 24998 24327 25050
rect 24165 24996 24189 24998
rect 24245 24996 24269 24998
rect 24325 24996 24349 24998
rect 24109 24976 24405 24996
rect 19478 24508 19774 24528
rect 19534 24506 19558 24508
rect 19614 24506 19638 24508
rect 19694 24506 19718 24508
rect 19556 24454 19558 24506
rect 19620 24454 19632 24506
rect 19694 24454 19696 24506
rect 19534 24452 19558 24454
rect 19614 24452 19638 24454
rect 19694 24452 19718 24454
rect 19478 24432 19774 24452
rect 14848 23964 15144 23984
rect 14904 23962 14928 23964
rect 14984 23962 15008 23964
rect 15064 23962 15088 23964
rect 14926 23910 14928 23962
rect 14990 23910 15002 23962
rect 15064 23910 15066 23962
rect 14904 23908 14928 23910
rect 14984 23908 15008 23910
rect 15064 23908 15088 23910
rect 14848 23888 15144 23908
rect 24109 23964 24405 23984
rect 24165 23962 24189 23964
rect 24245 23962 24269 23964
rect 24325 23962 24349 23964
rect 24187 23910 24189 23962
rect 24251 23910 24263 23962
rect 24325 23910 24327 23962
rect 24165 23908 24189 23910
rect 24245 23908 24269 23910
rect 24325 23908 24349 23910
rect 24109 23888 24405 23908
rect 19478 23420 19774 23440
rect 19534 23418 19558 23420
rect 19614 23418 19638 23420
rect 19694 23418 19718 23420
rect 19556 23366 19558 23418
rect 19620 23366 19632 23418
rect 19694 23366 19696 23418
rect 19534 23364 19558 23366
rect 19614 23364 19638 23366
rect 19694 23364 19718 23366
rect 19478 23344 19774 23364
rect 14848 22876 15144 22896
rect 14904 22874 14928 22876
rect 14984 22874 15008 22876
rect 15064 22874 15088 22876
rect 14926 22822 14928 22874
rect 14990 22822 15002 22874
rect 15064 22822 15066 22874
rect 14904 22820 14928 22822
rect 14984 22820 15008 22822
rect 15064 22820 15088 22822
rect 14848 22800 15144 22820
rect 24109 22876 24405 22896
rect 24165 22874 24189 22876
rect 24245 22874 24269 22876
rect 24325 22874 24349 22876
rect 24187 22822 24189 22874
rect 24251 22822 24263 22874
rect 24325 22822 24327 22874
rect 24165 22820 24189 22822
rect 24245 22820 24269 22822
rect 24325 22820 24349 22822
rect 24109 22800 24405 22820
rect 19478 22332 19774 22352
rect 19534 22330 19558 22332
rect 19614 22330 19638 22332
rect 19694 22330 19718 22332
rect 19556 22278 19558 22330
rect 19620 22278 19632 22330
rect 19694 22278 19696 22330
rect 19534 22276 19558 22278
rect 19614 22276 19638 22278
rect 19694 22276 19718 22278
rect 19478 22256 19774 22276
rect 14848 21788 15144 21808
rect 14904 21786 14928 21788
rect 14984 21786 15008 21788
rect 15064 21786 15088 21788
rect 14926 21734 14928 21786
rect 14990 21734 15002 21786
rect 15064 21734 15066 21786
rect 14904 21732 14928 21734
rect 14984 21732 15008 21734
rect 15064 21732 15088 21734
rect 14848 21712 15144 21732
rect 24109 21788 24405 21808
rect 24165 21786 24189 21788
rect 24245 21786 24269 21788
rect 24325 21786 24349 21788
rect 24187 21734 24189 21786
rect 24251 21734 24263 21786
rect 24325 21734 24327 21786
rect 24165 21732 24189 21734
rect 24245 21732 24269 21734
rect 24325 21732 24349 21734
rect 24109 21712 24405 21732
rect 19478 21244 19774 21264
rect 19534 21242 19558 21244
rect 19614 21242 19638 21244
rect 19694 21242 19718 21244
rect 19556 21190 19558 21242
rect 19620 21190 19632 21242
rect 19694 21190 19696 21242
rect 19534 21188 19558 21190
rect 19614 21188 19638 21190
rect 19694 21188 19718 21190
rect 19478 21168 19774 21188
rect 14848 20700 15144 20720
rect 14904 20698 14928 20700
rect 14984 20698 15008 20700
rect 15064 20698 15088 20700
rect 14926 20646 14928 20698
rect 14990 20646 15002 20698
rect 15064 20646 15066 20698
rect 14904 20644 14928 20646
rect 14984 20644 15008 20646
rect 15064 20644 15088 20646
rect 14848 20624 15144 20644
rect 24109 20700 24405 20720
rect 24165 20698 24189 20700
rect 24245 20698 24269 20700
rect 24325 20698 24349 20700
rect 24187 20646 24189 20698
rect 24251 20646 24263 20698
rect 24325 20646 24327 20698
rect 24165 20644 24189 20646
rect 24245 20644 24269 20646
rect 24325 20644 24349 20646
rect 24109 20624 24405 20644
rect 19478 20156 19774 20176
rect 19534 20154 19558 20156
rect 19614 20154 19638 20156
rect 19694 20154 19718 20156
rect 19556 20102 19558 20154
rect 19620 20102 19632 20154
rect 19694 20102 19696 20154
rect 19534 20100 19558 20102
rect 19614 20100 19638 20102
rect 19694 20100 19718 20102
rect 19478 20080 19774 20100
rect 14848 19612 15144 19632
rect 14904 19610 14928 19612
rect 14984 19610 15008 19612
rect 15064 19610 15088 19612
rect 14926 19558 14928 19610
rect 14990 19558 15002 19610
rect 15064 19558 15066 19610
rect 14904 19556 14928 19558
rect 14984 19556 15008 19558
rect 15064 19556 15088 19558
rect 14848 19536 15144 19556
rect 24109 19612 24405 19632
rect 24165 19610 24189 19612
rect 24245 19610 24269 19612
rect 24325 19610 24349 19612
rect 24187 19558 24189 19610
rect 24251 19558 24263 19610
rect 24325 19558 24327 19610
rect 24165 19556 24189 19558
rect 24245 19556 24269 19558
rect 24325 19556 24349 19558
rect 24109 19536 24405 19556
rect 19478 19068 19774 19088
rect 19534 19066 19558 19068
rect 19614 19066 19638 19068
rect 19694 19066 19718 19068
rect 19556 19014 19558 19066
rect 19620 19014 19632 19066
rect 19694 19014 19696 19066
rect 19534 19012 19558 19014
rect 19614 19012 19638 19014
rect 19694 19012 19718 19014
rect 19478 18992 19774 19012
rect 14848 18524 15144 18544
rect 14904 18522 14928 18524
rect 14984 18522 15008 18524
rect 15064 18522 15088 18524
rect 14926 18470 14928 18522
rect 14990 18470 15002 18522
rect 15064 18470 15066 18522
rect 14904 18468 14928 18470
rect 14984 18468 15008 18470
rect 15064 18468 15088 18470
rect 14848 18448 15144 18468
rect 24109 18524 24405 18544
rect 24165 18522 24189 18524
rect 24245 18522 24269 18524
rect 24325 18522 24349 18524
rect 24187 18470 24189 18522
rect 24251 18470 24263 18522
rect 24325 18470 24327 18522
rect 24165 18468 24189 18470
rect 24245 18468 24269 18470
rect 24325 18468 24349 18470
rect 24109 18448 24405 18468
rect 19478 17980 19774 18000
rect 19534 17978 19558 17980
rect 19614 17978 19638 17980
rect 19694 17978 19718 17980
rect 19556 17926 19558 17978
rect 19620 17926 19632 17978
rect 19694 17926 19696 17978
rect 19534 17924 19558 17926
rect 19614 17924 19638 17926
rect 19694 17924 19718 17926
rect 19478 17904 19774 17924
rect 14848 17436 15144 17456
rect 14904 17434 14928 17436
rect 14984 17434 15008 17436
rect 15064 17434 15088 17436
rect 14926 17382 14928 17434
rect 14990 17382 15002 17434
rect 15064 17382 15066 17434
rect 14904 17380 14928 17382
rect 14984 17380 15008 17382
rect 15064 17380 15088 17382
rect 14848 17360 15144 17380
rect 24109 17436 24405 17456
rect 24165 17434 24189 17436
rect 24245 17434 24269 17436
rect 24325 17434 24349 17436
rect 24187 17382 24189 17434
rect 24251 17382 24263 17434
rect 24325 17382 24327 17434
rect 24165 17380 24189 17382
rect 24245 17380 24269 17382
rect 24325 17380 24349 17382
rect 24109 17360 24405 17380
rect 28170 17096 28226 17105
rect 27988 17060 28040 17066
rect 28170 17031 28172 17040
rect 27988 17002 28040 17008
rect 28224 17031 28226 17040
rect 28172 17002 28224 17008
rect 19478 16892 19774 16912
rect 19534 16890 19558 16892
rect 19614 16890 19638 16892
rect 19694 16890 19718 16892
rect 19556 16838 19558 16890
rect 19620 16838 19632 16890
rect 19694 16838 19696 16890
rect 19534 16836 19558 16838
rect 19614 16836 19638 16838
rect 19694 16836 19718 16838
rect 19478 16816 19774 16836
rect 14848 16348 15144 16368
rect 14904 16346 14928 16348
rect 14984 16346 15008 16348
rect 15064 16346 15088 16348
rect 14926 16294 14928 16346
rect 14990 16294 15002 16346
rect 15064 16294 15066 16346
rect 14904 16292 14928 16294
rect 14984 16292 15008 16294
rect 15064 16292 15088 16294
rect 14848 16272 15144 16292
rect 24109 16348 24405 16368
rect 24165 16346 24189 16348
rect 24245 16346 24269 16348
rect 24325 16346 24349 16348
rect 24187 16294 24189 16346
rect 24251 16294 24263 16346
rect 24325 16294 24327 16346
rect 24165 16292 24189 16294
rect 24245 16292 24269 16294
rect 24325 16292 24349 16294
rect 24109 16272 24405 16292
rect 19478 15804 19774 15824
rect 19534 15802 19558 15804
rect 19614 15802 19638 15804
rect 19694 15802 19718 15804
rect 19556 15750 19558 15802
rect 19620 15750 19632 15802
rect 19694 15750 19696 15802
rect 19534 15748 19558 15750
rect 19614 15748 19638 15750
rect 19694 15748 19718 15750
rect 19478 15728 19774 15748
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13832 14958 13860 15302
rect 14848 15260 15144 15280
rect 14904 15258 14928 15260
rect 14984 15258 15008 15260
rect 15064 15258 15088 15260
rect 14926 15206 14928 15258
rect 14990 15206 15002 15258
rect 15064 15206 15066 15258
rect 14904 15204 14928 15206
rect 14984 15204 15008 15206
rect 15064 15204 15088 15206
rect 14848 15184 15144 15204
rect 24109 15260 24405 15280
rect 24165 15258 24189 15260
rect 24245 15258 24269 15260
rect 24325 15258 24349 15260
rect 24187 15206 24189 15258
rect 24251 15206 24263 15258
rect 24325 15206 24327 15258
rect 24165 15204 24189 15206
rect 24245 15204 24269 15206
rect 24325 15204 24349 15206
rect 24109 15184 24405 15204
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 10217 14716 10513 14736
rect 10273 14714 10297 14716
rect 10353 14714 10377 14716
rect 10433 14714 10457 14716
rect 10295 14662 10297 14714
rect 10359 14662 10371 14714
rect 10433 14662 10435 14714
rect 10273 14660 10297 14662
rect 10353 14660 10377 14662
rect 10433 14660 10457 14662
rect 10217 14640 10513 14660
rect 12268 14482 12296 14894
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12820 14482 12848 14758
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12084 14006 12112 14350
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 10217 13628 10513 13648
rect 10273 13626 10297 13628
rect 10353 13626 10377 13628
rect 10433 13626 10457 13628
rect 10295 13574 10297 13626
rect 10359 13574 10371 13626
rect 10433 13574 10435 13626
rect 10273 13572 10297 13574
rect 10353 13572 10377 13574
rect 10433 13572 10457 13574
rect 10217 13552 10513 13572
rect 12084 13326 12112 13942
rect 12164 13728 12216 13734
rect 12164 13670 12216 13676
rect 12176 13394 12204 13670
rect 12268 13530 12296 14418
rect 12912 13802 12940 14894
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 12900 13796 12952 13802
rect 12900 13738 12952 13744
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12912 13394 12940 13738
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 13096 13326 13124 14282
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 5586 13084 5882 13104
rect 5642 13082 5666 13084
rect 5722 13082 5746 13084
rect 5802 13082 5826 13084
rect 5664 13030 5666 13082
rect 5728 13030 5740 13082
rect 5802 13030 5804 13082
rect 5642 13028 5666 13030
rect 5722 13028 5746 13030
rect 5802 13028 5826 13030
rect 5586 13008 5882 13028
rect 13096 12986 13124 13262
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 5586 11996 5882 12016
rect 5642 11994 5666 11996
rect 5722 11994 5746 11996
rect 5802 11994 5826 11996
rect 5664 11942 5666 11994
rect 5728 11942 5740 11994
rect 5802 11942 5804 11994
rect 5642 11940 5666 11942
rect 5722 11940 5746 11942
rect 5802 11940 5826 11942
rect 5586 11920 5882 11940
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 11014 9720 11562
rect 9784 11218 9812 12174
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 5586 10908 5882 10928
rect 5642 10906 5666 10908
rect 5722 10906 5746 10908
rect 5802 10906 5826 10908
rect 5664 10854 5666 10906
rect 5728 10854 5740 10906
rect 5802 10854 5804 10906
rect 5642 10852 5666 10854
rect 5722 10852 5746 10854
rect 5802 10852 5826 10854
rect 5586 10832 5882 10852
rect 9692 10606 9720 10950
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9784 10062 9812 11154
rect 9968 10810 9996 12718
rect 10217 12540 10513 12560
rect 10273 12538 10297 12540
rect 10353 12538 10377 12540
rect 10433 12538 10457 12540
rect 10295 12486 10297 12538
rect 10359 12486 10371 12538
rect 10433 12486 10435 12538
rect 10273 12484 10297 12486
rect 10353 12484 10377 12486
rect 10433 12484 10457 12486
rect 10217 12464 10513 12484
rect 10980 11694 11008 12718
rect 12176 12374 12204 12718
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10217 11452 10513 11472
rect 10273 11450 10297 11452
rect 10353 11450 10377 11452
rect 10433 11450 10457 11452
rect 10295 11398 10297 11450
rect 10359 11398 10371 11450
rect 10433 11398 10435 11450
rect 10273 11396 10297 11398
rect 10353 11396 10377 11398
rect 10433 11396 10457 11398
rect 10217 11376 10513 11396
rect 10704 11286 10732 11494
rect 10692 11280 10744 11286
rect 10888 11268 10916 11630
rect 10968 11280 11020 11286
rect 10888 11240 10968 11268
rect 10692 11222 10744 11228
rect 10968 11222 11020 11228
rect 10980 10810 11008 11222
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11072 10742 11100 11766
rect 11532 11354 11560 12242
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 11532 10606 11560 11290
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11992 11098 12020 11154
rect 11900 11070 12020 11098
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 10600 10532 10652 10538
rect 10600 10474 10652 10480
rect 10217 10364 10513 10384
rect 10273 10362 10297 10364
rect 10353 10362 10377 10364
rect 10433 10362 10457 10364
rect 10295 10310 10297 10362
rect 10359 10310 10371 10362
rect 10433 10310 10435 10362
rect 10273 10308 10297 10310
rect 10353 10308 10377 10310
rect 10433 10308 10457 10310
rect 10217 10288 10513 10308
rect 10612 10266 10640 10474
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10600 10260 10652 10266
rect 10600 10202 10652 10208
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 5586 9820 5882 9840
rect 5642 9818 5666 9820
rect 5722 9818 5746 9820
rect 5802 9818 5826 9820
rect 5664 9766 5666 9818
rect 5728 9766 5740 9818
rect 5802 9766 5804 9818
rect 5642 9764 5666 9766
rect 5722 9764 5746 9766
rect 5802 9764 5826 9766
rect 5586 9744 5882 9764
rect 9784 9586 9812 9998
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 10152 9178 10180 10066
rect 10217 9276 10513 9296
rect 10273 9274 10297 9276
rect 10353 9274 10377 9276
rect 10433 9274 10457 9276
rect 10295 9222 10297 9274
rect 10359 9222 10371 9274
rect 10433 9222 10435 9274
rect 10273 9220 10297 9222
rect 10353 9220 10377 9222
rect 10433 9220 10457 9222
rect 10217 9200 10513 9220
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10612 9042 10640 10202
rect 10980 10198 11008 10406
rect 10968 10192 11020 10198
rect 10968 10134 11020 10140
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 5586 8732 5882 8752
rect 5642 8730 5666 8732
rect 5722 8730 5746 8732
rect 5802 8730 5826 8732
rect 5664 8678 5666 8730
rect 5728 8678 5740 8730
rect 5802 8678 5804 8730
rect 5642 8676 5666 8678
rect 5722 8676 5746 8678
rect 5802 8676 5826 8678
rect 5586 8656 5882 8676
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 5586 7644 5882 7664
rect 5642 7642 5666 7644
rect 5722 7642 5746 7644
rect 5802 7642 5826 7644
rect 5664 7590 5666 7642
rect 5728 7590 5740 7642
rect 5802 7590 5804 7642
rect 5642 7588 5666 7590
rect 5722 7588 5746 7590
rect 5802 7588 5826 7590
rect 5586 7568 5882 7588
rect 9784 7546 9812 7822
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 5586 6556 5882 6576
rect 5642 6554 5666 6556
rect 5722 6554 5746 6556
rect 5802 6554 5826 6556
rect 5664 6502 5666 6554
rect 5728 6502 5740 6554
rect 5802 6502 5804 6554
rect 5642 6500 5666 6502
rect 5722 6500 5746 6502
rect 5802 6500 5826 6502
rect 5586 6480 5882 6500
rect 10152 6254 10180 8842
rect 10888 8634 10916 9386
rect 10980 9178 11008 10134
rect 11900 9926 11928 11070
rect 12268 10810 12296 11630
rect 12452 11286 12480 12038
rect 12440 11280 12492 11286
rect 12440 11222 12492 11228
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12176 10130 12204 10406
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 11440 9042 11468 9862
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11532 9178 11560 9522
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11532 8838 11560 9114
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11532 8634 11560 8774
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 10217 8188 10513 8208
rect 10273 8186 10297 8188
rect 10353 8186 10377 8188
rect 10433 8186 10457 8188
rect 10295 8134 10297 8186
rect 10359 8134 10371 8186
rect 10433 8134 10435 8186
rect 10273 8132 10297 8134
rect 10353 8132 10377 8134
rect 10433 8132 10457 8134
rect 10217 8112 10513 8132
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 10612 7274 10640 7822
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7342 10916 7686
rect 10876 7336 10928 7342
rect 11060 7336 11112 7342
rect 10876 7278 10928 7284
rect 10980 7284 11060 7290
rect 10980 7278 11112 7284
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10980 7262 11100 7278
rect 10217 7100 10513 7120
rect 10273 7098 10297 7100
rect 10353 7098 10377 7100
rect 10433 7098 10457 7100
rect 10295 7046 10297 7098
rect 10359 7046 10371 7098
rect 10433 7046 10435 7098
rect 10273 7044 10297 7046
rect 10353 7044 10377 7046
rect 10433 7044 10457 7046
rect 10217 7024 10513 7044
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10217 6012 10513 6032
rect 10273 6010 10297 6012
rect 10353 6010 10377 6012
rect 10433 6010 10457 6012
rect 10295 5958 10297 6010
rect 10359 5958 10371 6010
rect 10433 5958 10435 6010
rect 10273 5956 10297 5958
rect 10353 5956 10377 5958
rect 10433 5956 10457 5958
rect 10217 5936 10513 5956
rect 10612 5846 10640 7210
rect 10980 6866 11008 7262
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10704 6118 10732 6802
rect 11716 6662 11744 7822
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11072 6186 11100 6598
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 5586 5468 5882 5488
rect 5642 5466 5666 5468
rect 5722 5466 5746 5468
rect 5802 5466 5826 5468
rect 5664 5414 5666 5466
rect 5728 5414 5740 5466
rect 5802 5414 5804 5466
rect 5642 5412 5666 5414
rect 5722 5412 5746 5414
rect 5802 5412 5826 5414
rect 5586 5392 5882 5412
rect 10060 4690 10088 5646
rect 10217 4924 10513 4944
rect 10273 4922 10297 4924
rect 10353 4922 10377 4924
rect 10433 4922 10457 4924
rect 10295 4870 10297 4922
rect 10359 4870 10371 4922
rect 10433 4870 10435 4922
rect 10273 4868 10297 4870
rect 10353 4868 10377 4870
rect 10433 4868 10457 4870
rect 10217 4848 10513 4868
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10600 4684 10652 4690
rect 10704 4672 10732 6054
rect 11532 5846 11560 6190
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 11072 4758 11100 4966
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 10652 4644 10732 4672
rect 10600 4626 10652 4632
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 5586 4380 5882 4400
rect 5642 4378 5666 4380
rect 5722 4378 5746 4380
rect 5802 4378 5826 4380
rect 5664 4326 5666 4378
rect 5728 4326 5740 4378
rect 5802 4326 5804 4378
rect 5642 4324 5666 4326
rect 5722 4324 5746 4326
rect 5802 4324 5826 4326
rect 5586 4304 5882 4324
rect 9968 3670 9996 4422
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10217 3836 10513 3856
rect 10273 3834 10297 3836
rect 10353 3834 10377 3836
rect 10433 3834 10457 3836
rect 10295 3782 10297 3834
rect 10359 3782 10371 3834
rect 10433 3782 10435 3834
rect 10273 3780 10297 3782
rect 10353 3780 10377 3782
rect 10433 3780 10457 3782
rect 10217 3760 10513 3780
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 5586 3292 5882 3312
rect 5642 3290 5666 3292
rect 5722 3290 5746 3292
rect 5802 3290 5826 3292
rect 5664 3238 5666 3290
rect 5728 3238 5740 3290
rect 5802 3238 5804 3290
rect 5642 3236 5666 3238
rect 5722 3236 5746 3238
rect 5802 3236 5826 3238
rect 5586 3216 5882 3236
rect 10217 2748 10513 2768
rect 10273 2746 10297 2748
rect 10353 2746 10377 2748
rect 10433 2746 10457 2748
rect 10295 2694 10297 2746
rect 10359 2694 10371 2746
rect 10433 2694 10435 2746
rect 10273 2692 10297 2694
rect 10353 2692 10377 2694
rect 10433 2692 10457 2694
rect 10217 2672 10513 2692
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 480 2508 532 2514
rect 480 2450 532 2456
rect 492 800 520 2450
rect 5586 2204 5882 2224
rect 5642 2202 5666 2204
rect 5722 2202 5746 2204
rect 5802 2202 5826 2204
rect 5664 2150 5666 2202
rect 5728 2150 5740 2202
rect 5802 2150 5804 2202
rect 5642 2148 5666 2150
rect 5722 2148 5746 2150
rect 5802 2148 5826 2150
rect 5586 2128 5882 2148
rect 10612 800 10640 3946
rect 10704 3602 10732 4644
rect 11164 4078 11192 5714
rect 11532 5166 11560 5782
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11808 4010 11836 8978
rect 11900 8430 11928 9862
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11888 6724 11940 6730
rect 11888 6666 11940 6672
rect 11900 6458 11928 6666
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11992 5778 12020 10066
rect 12176 9722 12204 10066
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12084 8430 12112 9386
rect 12268 8430 12296 9454
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12360 8090 12388 11018
rect 12544 10810 12572 12582
rect 12636 12442 12664 12650
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12912 11898 12940 12174
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 12728 11354 12756 11698
rect 13004 11354 13032 12174
rect 13096 11694 13124 12922
rect 13188 12306 13216 13806
rect 13360 12436 13412 12442
rect 13360 12378 13412 12384
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 13280 11898 13308 12106
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13372 11778 13400 12378
rect 13464 12374 13492 13806
rect 13556 12434 13584 14214
rect 13740 12442 13768 14758
rect 13832 14482 13860 14894
rect 19478 14716 19774 14736
rect 19534 14714 19558 14716
rect 19614 14714 19638 14716
rect 19694 14714 19718 14716
rect 19556 14662 19558 14714
rect 19620 14662 19632 14714
rect 19694 14662 19696 14714
rect 19534 14660 19558 14662
rect 19614 14660 19638 14662
rect 19694 14660 19718 14662
rect 19478 14640 19774 14660
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 14848 14172 15144 14192
rect 14904 14170 14928 14172
rect 14984 14170 15008 14172
rect 15064 14170 15088 14172
rect 14926 14118 14928 14170
rect 14990 14118 15002 14170
rect 15064 14118 15066 14170
rect 14904 14116 14928 14118
rect 14984 14116 15008 14118
rect 15064 14116 15088 14118
rect 14848 14096 15144 14116
rect 24109 14172 24405 14192
rect 24165 14170 24189 14172
rect 24245 14170 24269 14172
rect 24325 14170 24349 14172
rect 24187 14118 24189 14170
rect 24251 14118 24263 14170
rect 24325 14118 24327 14170
rect 24165 14116 24189 14118
rect 24245 14116 24269 14118
rect 24325 14116 24349 14118
rect 24109 14096 24405 14116
rect 28000 13870 28028 17002
rect 27988 13864 28040 13870
rect 27988 13806 28040 13812
rect 14372 13796 14424 13802
rect 14372 13738 14424 13744
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 12782 14044 13126
rect 14384 12986 14412 13738
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 13394 15332 13670
rect 19478 13628 19774 13648
rect 19534 13626 19558 13628
rect 19614 13626 19638 13628
rect 19694 13626 19718 13628
rect 19556 13574 19558 13626
rect 19620 13574 19632 13626
rect 19694 13574 19696 13626
rect 19534 13572 19558 13574
rect 19614 13572 19638 13574
rect 19694 13572 19718 13574
rect 19478 13552 19774 13572
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 14848 13084 15144 13104
rect 14904 13082 14928 13084
rect 14984 13082 15008 13084
rect 15064 13082 15088 13084
rect 14926 13030 14928 13082
rect 14990 13030 15002 13082
rect 15064 13030 15066 13082
rect 14904 13028 14928 13030
rect 14984 13028 15008 13030
rect 15064 13028 15088 13030
rect 14848 13008 15144 13028
rect 24109 13084 24405 13104
rect 24165 13082 24189 13084
rect 24245 13082 24269 13084
rect 24325 13082 24349 13084
rect 24187 13030 24189 13082
rect 24251 13030 24263 13082
rect 24325 13030 24327 13082
rect 24165 13028 24189 13030
rect 24245 13028 24269 13030
rect 24325 13028 24349 13030
rect 24109 13008 24405 13028
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14556 12708 14608 12714
rect 14556 12650 14608 12656
rect 13728 12436 13780 12442
rect 13556 12406 13676 12434
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13464 12102 13492 12310
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13648 11778 13676 12406
rect 14568 12434 14596 12650
rect 19478 12540 19774 12560
rect 19534 12538 19558 12540
rect 19614 12538 19638 12540
rect 19694 12538 19718 12540
rect 19556 12486 19558 12538
rect 19620 12486 19632 12538
rect 19694 12486 19696 12538
rect 19534 12484 19558 12486
rect 19614 12484 19638 12486
rect 19694 12484 19718 12486
rect 19478 12464 19774 12484
rect 13728 12378 13780 12384
rect 14476 12406 14596 12434
rect 14476 12374 14504 12406
rect 14464 12368 14516 12374
rect 14464 12310 14516 12316
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13280 11750 13400 11778
rect 13464 11750 13676 11778
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12164 8016 12216 8022
rect 12164 7958 12216 7964
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12084 6934 12112 7686
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 12084 6254 12112 6870
rect 12176 6866 12204 7958
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12268 7546 12296 7754
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 12176 5914 12204 6802
rect 12360 6798 12388 7686
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12452 6458 12480 6802
rect 12544 6662 12572 7890
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12728 6798 12756 7142
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12728 6254 12756 6734
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 12268 5234 12296 6054
rect 12360 5846 12388 6122
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 12360 5370 12388 5782
rect 12820 5370 12848 7890
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12912 5778 12940 7210
rect 13280 6866 13308 11750
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13372 11014 13400 11630
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13372 10810 13400 10950
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13464 7936 13492 11750
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13556 10674 13584 11086
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13464 7908 13584 7936
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 13464 7342 13492 7754
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13280 6186 13308 6802
rect 13372 6662 13400 7210
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 6254 13400 6598
rect 13464 6458 13492 7278
rect 13556 6866 13584 7908
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13268 6180 13320 6186
rect 13268 6122 13320 6128
rect 13372 5846 13400 6190
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 12176 4078 12204 4694
rect 12164 4072 12216 4078
rect 12164 4014 12216 4020
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 12268 3194 12296 5170
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12360 4758 12388 5102
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 12544 4690 12572 5170
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12636 4690 12664 5102
rect 12728 4826 12756 5102
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12360 3942 12388 4558
rect 12544 4282 12572 4626
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 12544 2990 12572 4218
rect 12636 4146 12664 4626
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12636 3058 12664 4082
rect 12820 4010 12848 4150
rect 12912 4078 12940 4762
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12912 3398 12940 4014
rect 13004 3942 13032 5714
rect 13556 5574 13584 6802
rect 13648 6730 13676 11630
rect 13740 8906 13768 12242
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13832 10810 13860 11154
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13832 10538 13860 10746
rect 13820 10532 13872 10538
rect 13820 10474 13872 10480
rect 14108 10470 14136 11834
rect 14476 11626 14504 12310
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14292 10810 14320 11494
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14188 10600 14240 10606
rect 14240 10548 14412 10554
rect 14188 10542 14412 10548
rect 14200 10538 14412 10542
rect 14200 10532 14424 10538
rect 14200 10526 14372 10532
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13832 9518 13860 9930
rect 13924 9586 13952 10406
rect 14200 10130 14228 10406
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14292 9722 14320 10526
rect 14372 10474 14424 10480
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 14476 9450 14504 11562
rect 14568 11218 14596 12038
rect 14660 11694 14688 12038
rect 14848 11996 15144 12016
rect 14904 11994 14928 11996
rect 14984 11994 15008 11996
rect 15064 11994 15088 11996
rect 14926 11942 14928 11994
rect 14990 11942 15002 11994
rect 15064 11942 15066 11994
rect 14904 11940 14928 11942
rect 14984 11940 15008 11942
rect 15064 11940 15088 11942
rect 14848 11920 15144 11940
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14660 11286 14688 11630
rect 14648 11280 14700 11286
rect 14648 11222 14700 11228
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14568 10690 14596 11154
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 15120 11098 15148 11698
rect 15580 11558 15608 12174
rect 24109 11996 24405 12016
rect 24165 11994 24189 11996
rect 24245 11994 24269 11996
rect 24325 11994 24349 11996
rect 24187 11942 24189 11994
rect 24251 11942 24263 11994
rect 24325 11942 24327 11994
rect 24165 11940 24189 11942
rect 24245 11940 24269 11942
rect 24325 11940 24349 11942
rect 24109 11920 24405 11940
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 14660 10810 14688 11086
rect 15120 11070 15240 11098
rect 14848 10908 15144 10928
rect 14904 10906 14928 10908
rect 14984 10906 15008 10908
rect 15064 10906 15088 10908
rect 14926 10854 14928 10906
rect 14990 10854 15002 10906
rect 15064 10854 15066 10906
rect 14904 10852 14928 10854
rect 14984 10852 15008 10854
rect 15064 10852 15088 10854
rect 14848 10832 15144 10852
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 15212 10724 15240 11070
rect 15384 10736 15436 10742
rect 14752 10696 15384 10724
rect 14568 10662 14688 10690
rect 14660 10062 14688 10662
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13832 7410 13860 7822
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13832 6254 13860 7346
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13832 5250 13860 5850
rect 13924 5778 13952 7346
rect 14476 7206 14504 9386
rect 14660 9042 14688 9998
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14568 7274 14596 8366
rect 14752 8022 14780 10696
rect 15384 10678 15436 10684
rect 15580 10538 15608 11494
rect 16132 11354 16160 11630
rect 19478 11452 19774 11472
rect 19534 11450 19558 11452
rect 19614 11450 19638 11452
rect 19694 11450 19718 11452
rect 19556 11398 19558 11450
rect 19620 11398 19632 11450
rect 19694 11398 19696 11450
rect 19534 11396 19558 11398
rect 19614 11396 19638 11398
rect 19694 11396 19718 11398
rect 19478 11376 19774 11396
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 24109 10908 24405 10928
rect 24165 10906 24189 10908
rect 24245 10906 24269 10908
rect 24325 10906 24349 10908
rect 24187 10854 24189 10906
rect 24251 10854 24263 10906
rect 24325 10854 24327 10906
rect 24165 10852 24189 10854
rect 24245 10852 24269 10854
rect 24325 10852 24349 10854
rect 24109 10832 24405 10852
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 16132 10266 16160 10610
rect 19478 10364 19774 10384
rect 19534 10362 19558 10364
rect 19614 10362 19638 10364
rect 19694 10362 19718 10364
rect 19556 10310 19558 10362
rect 19620 10310 19632 10362
rect 19694 10310 19696 10362
rect 19534 10308 19558 10310
rect 19614 10308 19638 10310
rect 19694 10308 19718 10310
rect 19478 10288 19774 10308
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 14848 9820 15144 9840
rect 14904 9818 14928 9820
rect 14984 9818 15008 9820
rect 15064 9818 15088 9820
rect 14926 9766 14928 9818
rect 14990 9766 15002 9818
rect 15064 9766 15066 9818
rect 14904 9764 14928 9766
rect 14984 9764 15008 9766
rect 15064 9764 15088 9766
rect 14848 9744 15144 9764
rect 24109 9820 24405 9840
rect 24165 9818 24189 9820
rect 24245 9818 24269 9820
rect 24325 9818 24349 9820
rect 24187 9766 24189 9818
rect 24251 9766 24263 9818
rect 24325 9766 24327 9818
rect 24165 9764 24189 9766
rect 24245 9764 24269 9766
rect 24325 9764 24349 9766
rect 24109 9744 24405 9764
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 14848 8732 15144 8752
rect 14904 8730 14928 8732
rect 14984 8730 15008 8732
rect 15064 8730 15088 8732
rect 14926 8678 14928 8730
rect 14990 8678 15002 8730
rect 15064 8678 15066 8730
rect 14904 8676 14928 8678
rect 14984 8676 15008 8678
rect 15064 8676 15088 8678
rect 14848 8656 15144 8676
rect 15212 8430 15240 9454
rect 15304 8498 15332 9522
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16132 9110 16160 9318
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 16224 8922 16252 9386
rect 19478 9276 19774 9296
rect 19534 9274 19558 9276
rect 19614 9274 19638 9276
rect 19694 9274 19718 9276
rect 19556 9222 19558 9274
rect 19620 9222 19632 9274
rect 19694 9222 19696 9274
rect 19534 9220 19558 9222
rect 19614 9220 19638 9222
rect 19694 9220 19718 9222
rect 19478 9200 19774 9220
rect 16132 8894 16252 8922
rect 16132 8838 16160 8894
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 16132 8430 16160 8774
rect 24109 8732 24405 8752
rect 24165 8730 24189 8732
rect 24245 8730 24269 8732
rect 24325 8730 24349 8732
rect 24187 8678 24189 8730
rect 24251 8678 24263 8730
rect 24325 8678 24327 8730
rect 24165 8676 24189 8678
rect 24245 8676 24269 8678
rect 24325 8676 24349 8678
rect 24109 8656 24405 8676
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 19478 8188 19774 8208
rect 19534 8186 19558 8188
rect 19614 8186 19638 8188
rect 19694 8186 19718 8188
rect 19556 8134 19558 8186
rect 19620 8134 19632 8186
rect 19694 8134 19696 8186
rect 19534 8132 19558 8134
rect 19614 8132 19638 8134
rect 19694 8132 19718 8134
rect 19478 8112 19774 8132
rect 14740 8016 14792 8022
rect 14740 7958 14792 7964
rect 14752 7546 14780 7958
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 14848 7644 15144 7664
rect 14904 7642 14928 7644
rect 14984 7642 15008 7644
rect 15064 7642 15088 7644
rect 14926 7590 14928 7642
rect 14990 7590 15002 7642
rect 15064 7590 15066 7642
rect 14904 7588 14928 7590
rect 14984 7588 15008 7590
rect 15064 7588 15088 7590
rect 14848 7568 15144 7588
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15120 7342 15148 7414
rect 15396 7342 15424 7686
rect 24109 7644 24405 7664
rect 24165 7642 24189 7644
rect 24245 7642 24269 7644
rect 24325 7642 24349 7644
rect 24187 7590 24189 7642
rect 24251 7590 24263 7642
rect 24325 7590 24327 7642
rect 24165 7588 24189 7590
rect 24245 7588 24269 7590
rect 24325 7588 24349 7590
rect 24109 7568 24405 7588
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15028 6866 15056 7142
rect 19478 7100 19774 7120
rect 19534 7098 19558 7100
rect 19614 7098 19638 7100
rect 19694 7098 19718 7100
rect 19556 7046 19558 7098
rect 19620 7046 19632 7098
rect 19694 7046 19696 7098
rect 19534 7044 19558 7046
rect 19614 7044 19638 7046
rect 19694 7044 19718 7046
rect 19478 7024 19774 7044
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13648 5222 13860 5250
rect 13648 5166 13676 5222
rect 13636 5160 13688 5166
rect 13820 5160 13872 5166
rect 13636 5102 13688 5108
rect 13740 5120 13820 5148
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13268 4548 13320 4554
rect 13268 4490 13320 4496
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13280 3738 13308 4490
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 13280 2990 13308 3674
rect 13556 3602 13584 4966
rect 13740 4010 13768 5120
rect 13820 5102 13872 5108
rect 13924 4826 13952 5714
rect 14476 5642 14504 6598
rect 14752 5914 14780 6734
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 14848 6556 15144 6576
rect 14904 6554 14928 6556
rect 14984 6554 15008 6556
rect 15064 6554 15088 6556
rect 14926 6502 14928 6554
rect 14990 6502 15002 6554
rect 15064 6502 15066 6554
rect 14904 6500 14928 6502
rect 14984 6500 15008 6502
rect 15064 6500 15088 6502
rect 14848 6480 15144 6500
rect 15396 6254 15424 6598
rect 24109 6556 24405 6576
rect 24165 6554 24189 6556
rect 24245 6554 24269 6556
rect 24325 6554 24349 6556
rect 24187 6502 24189 6554
rect 24251 6502 24263 6554
rect 24325 6502 24327 6554
rect 24165 6500 24189 6502
rect 24245 6500 24269 6502
rect 24325 6500 24349 6502
rect 24109 6480 24405 6500
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 16396 6180 16448 6186
rect 16396 6122 16448 6128
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14936 5778 14964 6054
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 14016 4690 14044 5170
rect 14476 5166 14504 5578
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 14848 5468 15144 5488
rect 14904 5466 14928 5468
rect 14984 5466 15008 5468
rect 15064 5466 15088 5468
rect 14926 5414 14928 5466
rect 14990 5414 15002 5466
rect 15064 5414 15066 5466
rect 14904 5412 14928 5414
rect 14984 5412 15008 5414
rect 15064 5412 15088 5414
rect 14848 5392 15144 5412
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14384 4282 14412 4558
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13832 3602 13860 4014
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 14384 2990 14412 4218
rect 14752 3738 14780 4626
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 14848 4380 15144 4400
rect 14904 4378 14928 4380
rect 14984 4378 15008 4380
rect 15064 4378 15088 4380
rect 14926 4326 14928 4378
rect 14990 4326 15002 4378
rect 15064 4326 15066 4378
rect 14904 4324 14928 4326
rect 14984 4324 15008 4326
rect 15064 4324 15088 4326
rect 14848 4304 15144 4324
rect 15304 4078 15332 4422
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 15672 3534 15700 5510
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15856 3738 15884 4422
rect 15948 4282 15976 5102
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16224 4826 16252 4966
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16408 4622 16436 6122
rect 19478 6012 19774 6032
rect 19534 6010 19558 6012
rect 19614 6010 19638 6012
rect 19694 6010 19718 6012
rect 19556 5958 19558 6010
rect 19620 5958 19632 6010
rect 19694 5958 19696 6010
rect 19534 5956 19558 5958
rect 19614 5956 19638 5958
rect 19694 5956 19718 5958
rect 19478 5936 19774 5956
rect 24109 5468 24405 5488
rect 24165 5466 24189 5468
rect 24245 5466 24269 5468
rect 24325 5466 24349 5468
rect 24187 5414 24189 5466
rect 24251 5414 24263 5466
rect 24325 5414 24327 5466
rect 24165 5412 24189 5414
rect 24245 5412 24269 5414
rect 24325 5412 24349 5414
rect 24109 5392 24405 5412
rect 19478 4924 19774 4944
rect 19534 4922 19558 4924
rect 19614 4922 19638 4924
rect 19694 4922 19718 4924
rect 19556 4870 19558 4922
rect 19620 4870 19632 4922
rect 19694 4870 19696 4922
rect 19534 4868 19558 4870
rect 19614 4868 19638 4870
rect 19694 4868 19718 4870
rect 19478 4848 19774 4868
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 14848 3292 15144 3312
rect 14904 3290 14928 3292
rect 14984 3290 15008 3292
rect 15064 3290 15088 3292
rect 14926 3238 14928 3290
rect 14990 3238 15002 3290
rect 15064 3238 15066 3290
rect 14904 3236 14928 3238
rect 14984 3236 15008 3238
rect 15064 3236 15088 3238
rect 14848 3216 15144 3236
rect 17880 3194 17908 4626
rect 24109 4380 24405 4400
rect 24165 4378 24189 4380
rect 24245 4378 24269 4380
rect 24325 4378 24349 4380
rect 24187 4326 24189 4378
rect 24251 4326 24263 4378
rect 24325 4326 24327 4378
rect 24165 4324 24189 4326
rect 24245 4324 24269 4326
rect 24325 4324 24349 4326
rect 24109 4304 24405 4324
rect 19478 3836 19774 3856
rect 19534 3834 19558 3836
rect 19614 3834 19638 3836
rect 19694 3834 19718 3836
rect 19556 3782 19558 3834
rect 19620 3782 19632 3834
rect 19694 3782 19696 3834
rect 19534 3780 19558 3782
rect 19614 3780 19638 3782
rect 19694 3780 19718 3782
rect 19478 3760 19774 3780
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 24109 3292 24405 3312
rect 24165 3290 24189 3292
rect 24245 3290 24269 3292
rect 24325 3290 24349 3292
rect 24187 3238 24189 3290
rect 24251 3238 24263 3290
rect 24325 3238 24327 3290
rect 24165 3236 24189 3238
rect 24245 3236 24269 3238
rect 24325 3236 24349 3238
rect 24109 3216 24405 3236
rect 27908 3194 27936 3470
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 27896 3188 27948 3194
rect 27896 3130 27948 3136
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 27344 2984 27396 2990
rect 27344 2926 27396 2932
rect 19478 2748 19774 2768
rect 19534 2746 19558 2748
rect 19614 2746 19638 2748
rect 19694 2746 19718 2748
rect 19556 2694 19558 2746
rect 19620 2694 19632 2746
rect 19694 2694 19696 2746
rect 19534 2692 19558 2694
rect 19614 2692 19638 2694
rect 19694 2692 19718 2694
rect 19478 2672 19774 2692
rect 20732 2650 20760 2926
rect 27356 2650 27384 2926
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 27160 2508 27212 2514
rect 27160 2450 27212 2456
rect 14848 2204 15144 2224
rect 14904 2202 14928 2204
rect 14984 2202 15008 2204
rect 15064 2202 15088 2204
rect 14926 2150 14928 2202
rect 14990 2150 15002 2202
rect 15064 2150 15066 2202
rect 14904 2148 14928 2150
rect 14984 2148 15008 2150
rect 15064 2148 15088 2150
rect 14848 2128 15144 2148
rect 20732 800 20760 2450
rect 24109 2204 24405 2224
rect 24165 2202 24189 2204
rect 24245 2202 24269 2204
rect 24325 2202 24349 2204
rect 24187 2150 24189 2202
rect 24251 2150 24263 2202
rect 24325 2150 24327 2202
rect 24165 2148 24189 2150
rect 24245 2148 24269 2150
rect 24325 2148 24349 2150
rect 24109 2128 24405 2148
rect 27172 2145 27200 2450
rect 27158 2136 27214 2145
rect 27158 2071 27214 2080
rect 478 0 534 800
rect 10598 0 10654 800
rect 20718 0 20774 800
<< via2 >>
rect 1398 29960 1454 30016
rect 10217 29946 10273 29948
rect 10297 29946 10353 29948
rect 10377 29946 10433 29948
rect 10457 29946 10513 29948
rect 10217 29894 10243 29946
rect 10243 29894 10273 29946
rect 10297 29894 10307 29946
rect 10307 29894 10353 29946
rect 10377 29894 10423 29946
rect 10423 29894 10433 29946
rect 10457 29894 10487 29946
rect 10487 29894 10513 29946
rect 10217 29892 10273 29894
rect 10297 29892 10353 29894
rect 10377 29892 10433 29894
rect 10457 29892 10513 29894
rect 19478 29946 19534 29948
rect 19558 29946 19614 29948
rect 19638 29946 19694 29948
rect 19718 29946 19774 29948
rect 19478 29894 19504 29946
rect 19504 29894 19534 29946
rect 19558 29894 19568 29946
rect 19568 29894 19614 29946
rect 19638 29894 19684 29946
rect 19684 29894 19694 29946
rect 19718 29894 19748 29946
rect 19748 29894 19774 29946
rect 19478 29892 19534 29894
rect 19558 29892 19614 29894
rect 19638 29892 19694 29894
rect 19718 29892 19774 29894
rect 1398 15000 1454 15056
rect 5586 29402 5642 29404
rect 5666 29402 5722 29404
rect 5746 29402 5802 29404
rect 5826 29402 5882 29404
rect 5586 29350 5612 29402
rect 5612 29350 5642 29402
rect 5666 29350 5676 29402
rect 5676 29350 5722 29402
rect 5746 29350 5792 29402
rect 5792 29350 5802 29402
rect 5826 29350 5856 29402
rect 5856 29350 5882 29402
rect 5586 29348 5642 29350
rect 5666 29348 5722 29350
rect 5746 29348 5802 29350
rect 5826 29348 5882 29350
rect 5586 28314 5642 28316
rect 5666 28314 5722 28316
rect 5746 28314 5802 28316
rect 5826 28314 5882 28316
rect 5586 28262 5612 28314
rect 5612 28262 5642 28314
rect 5666 28262 5676 28314
rect 5676 28262 5722 28314
rect 5746 28262 5792 28314
rect 5792 28262 5802 28314
rect 5826 28262 5856 28314
rect 5856 28262 5882 28314
rect 5586 28260 5642 28262
rect 5666 28260 5722 28262
rect 5746 28260 5802 28262
rect 5826 28260 5882 28262
rect 5586 27226 5642 27228
rect 5666 27226 5722 27228
rect 5746 27226 5802 27228
rect 5826 27226 5882 27228
rect 5586 27174 5612 27226
rect 5612 27174 5642 27226
rect 5666 27174 5676 27226
rect 5676 27174 5722 27226
rect 5746 27174 5792 27226
rect 5792 27174 5802 27226
rect 5826 27174 5856 27226
rect 5856 27174 5882 27226
rect 5586 27172 5642 27174
rect 5666 27172 5722 27174
rect 5746 27172 5802 27174
rect 5826 27172 5882 27174
rect 5586 26138 5642 26140
rect 5666 26138 5722 26140
rect 5746 26138 5802 26140
rect 5826 26138 5882 26140
rect 5586 26086 5612 26138
rect 5612 26086 5642 26138
rect 5666 26086 5676 26138
rect 5676 26086 5722 26138
rect 5746 26086 5792 26138
rect 5792 26086 5802 26138
rect 5826 26086 5856 26138
rect 5856 26086 5882 26138
rect 5586 26084 5642 26086
rect 5666 26084 5722 26086
rect 5746 26084 5802 26086
rect 5826 26084 5882 26086
rect 5586 25050 5642 25052
rect 5666 25050 5722 25052
rect 5746 25050 5802 25052
rect 5826 25050 5882 25052
rect 5586 24998 5612 25050
rect 5612 24998 5642 25050
rect 5666 24998 5676 25050
rect 5676 24998 5722 25050
rect 5746 24998 5792 25050
rect 5792 24998 5802 25050
rect 5826 24998 5856 25050
rect 5856 24998 5882 25050
rect 5586 24996 5642 24998
rect 5666 24996 5722 24998
rect 5746 24996 5802 24998
rect 5826 24996 5882 24998
rect 5586 23962 5642 23964
rect 5666 23962 5722 23964
rect 5746 23962 5802 23964
rect 5826 23962 5882 23964
rect 5586 23910 5612 23962
rect 5612 23910 5642 23962
rect 5666 23910 5676 23962
rect 5676 23910 5722 23962
rect 5746 23910 5792 23962
rect 5792 23910 5802 23962
rect 5826 23910 5856 23962
rect 5856 23910 5882 23962
rect 5586 23908 5642 23910
rect 5666 23908 5722 23910
rect 5746 23908 5802 23910
rect 5826 23908 5882 23910
rect 5586 22874 5642 22876
rect 5666 22874 5722 22876
rect 5746 22874 5802 22876
rect 5826 22874 5882 22876
rect 5586 22822 5612 22874
rect 5612 22822 5642 22874
rect 5666 22822 5676 22874
rect 5676 22822 5722 22874
rect 5746 22822 5792 22874
rect 5792 22822 5802 22874
rect 5826 22822 5856 22874
rect 5856 22822 5882 22874
rect 5586 22820 5642 22822
rect 5666 22820 5722 22822
rect 5746 22820 5802 22822
rect 5826 22820 5882 22822
rect 5586 21786 5642 21788
rect 5666 21786 5722 21788
rect 5746 21786 5802 21788
rect 5826 21786 5882 21788
rect 5586 21734 5612 21786
rect 5612 21734 5642 21786
rect 5666 21734 5676 21786
rect 5676 21734 5722 21786
rect 5746 21734 5792 21786
rect 5792 21734 5802 21786
rect 5826 21734 5856 21786
rect 5856 21734 5882 21786
rect 5586 21732 5642 21734
rect 5666 21732 5722 21734
rect 5746 21732 5802 21734
rect 5826 21732 5882 21734
rect 5586 20698 5642 20700
rect 5666 20698 5722 20700
rect 5746 20698 5802 20700
rect 5826 20698 5882 20700
rect 5586 20646 5612 20698
rect 5612 20646 5642 20698
rect 5666 20646 5676 20698
rect 5676 20646 5722 20698
rect 5746 20646 5792 20698
rect 5792 20646 5802 20698
rect 5826 20646 5856 20698
rect 5856 20646 5882 20698
rect 5586 20644 5642 20646
rect 5666 20644 5722 20646
rect 5746 20644 5802 20646
rect 5826 20644 5882 20646
rect 5586 19610 5642 19612
rect 5666 19610 5722 19612
rect 5746 19610 5802 19612
rect 5826 19610 5882 19612
rect 5586 19558 5612 19610
rect 5612 19558 5642 19610
rect 5666 19558 5676 19610
rect 5676 19558 5722 19610
rect 5746 19558 5792 19610
rect 5792 19558 5802 19610
rect 5826 19558 5856 19610
rect 5856 19558 5882 19610
rect 5586 19556 5642 19558
rect 5666 19556 5722 19558
rect 5746 19556 5802 19558
rect 5826 19556 5882 19558
rect 5586 18522 5642 18524
rect 5666 18522 5722 18524
rect 5746 18522 5802 18524
rect 5826 18522 5882 18524
rect 5586 18470 5612 18522
rect 5612 18470 5642 18522
rect 5666 18470 5676 18522
rect 5676 18470 5722 18522
rect 5746 18470 5792 18522
rect 5792 18470 5802 18522
rect 5826 18470 5856 18522
rect 5856 18470 5882 18522
rect 5586 18468 5642 18470
rect 5666 18468 5722 18470
rect 5746 18468 5802 18470
rect 5826 18468 5882 18470
rect 5586 17434 5642 17436
rect 5666 17434 5722 17436
rect 5746 17434 5802 17436
rect 5826 17434 5882 17436
rect 5586 17382 5612 17434
rect 5612 17382 5642 17434
rect 5666 17382 5676 17434
rect 5676 17382 5722 17434
rect 5746 17382 5792 17434
rect 5792 17382 5802 17434
rect 5826 17382 5856 17434
rect 5856 17382 5882 17434
rect 5586 17380 5642 17382
rect 5666 17380 5722 17382
rect 5746 17380 5802 17382
rect 5826 17380 5882 17382
rect 5586 16346 5642 16348
rect 5666 16346 5722 16348
rect 5746 16346 5802 16348
rect 5826 16346 5882 16348
rect 5586 16294 5612 16346
rect 5612 16294 5642 16346
rect 5666 16294 5676 16346
rect 5676 16294 5722 16346
rect 5746 16294 5792 16346
rect 5792 16294 5802 16346
rect 5826 16294 5856 16346
rect 5856 16294 5882 16346
rect 5586 16292 5642 16294
rect 5666 16292 5722 16294
rect 5746 16292 5802 16294
rect 5826 16292 5882 16294
rect 5586 15258 5642 15260
rect 5666 15258 5722 15260
rect 5746 15258 5802 15260
rect 5826 15258 5882 15260
rect 5586 15206 5612 15258
rect 5612 15206 5642 15258
rect 5666 15206 5676 15258
rect 5676 15206 5722 15258
rect 5746 15206 5792 15258
rect 5792 15206 5802 15258
rect 5826 15206 5856 15258
rect 5856 15206 5882 15258
rect 5586 15204 5642 15206
rect 5666 15204 5722 15206
rect 5746 15204 5802 15206
rect 5826 15204 5882 15206
rect 5586 14170 5642 14172
rect 5666 14170 5722 14172
rect 5746 14170 5802 14172
rect 5826 14170 5882 14172
rect 5586 14118 5612 14170
rect 5612 14118 5642 14170
rect 5666 14118 5676 14170
rect 5676 14118 5722 14170
rect 5746 14118 5792 14170
rect 5792 14118 5802 14170
rect 5826 14118 5856 14170
rect 5856 14118 5882 14170
rect 5586 14116 5642 14118
rect 5666 14116 5722 14118
rect 5746 14116 5802 14118
rect 5826 14116 5882 14118
rect 10217 28858 10273 28860
rect 10297 28858 10353 28860
rect 10377 28858 10433 28860
rect 10457 28858 10513 28860
rect 10217 28806 10243 28858
rect 10243 28806 10273 28858
rect 10297 28806 10307 28858
rect 10307 28806 10353 28858
rect 10377 28806 10423 28858
rect 10423 28806 10433 28858
rect 10457 28806 10487 28858
rect 10487 28806 10513 28858
rect 10217 28804 10273 28806
rect 10297 28804 10353 28806
rect 10377 28804 10433 28806
rect 10457 28804 10513 28806
rect 10217 27770 10273 27772
rect 10297 27770 10353 27772
rect 10377 27770 10433 27772
rect 10457 27770 10513 27772
rect 10217 27718 10243 27770
rect 10243 27718 10273 27770
rect 10297 27718 10307 27770
rect 10307 27718 10353 27770
rect 10377 27718 10423 27770
rect 10423 27718 10433 27770
rect 10457 27718 10487 27770
rect 10487 27718 10513 27770
rect 10217 27716 10273 27718
rect 10297 27716 10353 27718
rect 10377 27716 10433 27718
rect 10457 27716 10513 27718
rect 10217 26682 10273 26684
rect 10297 26682 10353 26684
rect 10377 26682 10433 26684
rect 10457 26682 10513 26684
rect 10217 26630 10243 26682
rect 10243 26630 10273 26682
rect 10297 26630 10307 26682
rect 10307 26630 10353 26682
rect 10377 26630 10423 26682
rect 10423 26630 10433 26682
rect 10457 26630 10487 26682
rect 10487 26630 10513 26682
rect 10217 26628 10273 26630
rect 10297 26628 10353 26630
rect 10377 26628 10433 26630
rect 10457 26628 10513 26630
rect 10217 25594 10273 25596
rect 10297 25594 10353 25596
rect 10377 25594 10433 25596
rect 10457 25594 10513 25596
rect 10217 25542 10243 25594
rect 10243 25542 10273 25594
rect 10297 25542 10307 25594
rect 10307 25542 10353 25594
rect 10377 25542 10423 25594
rect 10423 25542 10433 25594
rect 10457 25542 10487 25594
rect 10487 25542 10513 25594
rect 10217 25540 10273 25542
rect 10297 25540 10353 25542
rect 10377 25540 10433 25542
rect 10457 25540 10513 25542
rect 10217 24506 10273 24508
rect 10297 24506 10353 24508
rect 10377 24506 10433 24508
rect 10457 24506 10513 24508
rect 10217 24454 10243 24506
rect 10243 24454 10273 24506
rect 10297 24454 10307 24506
rect 10307 24454 10353 24506
rect 10377 24454 10423 24506
rect 10423 24454 10433 24506
rect 10457 24454 10487 24506
rect 10487 24454 10513 24506
rect 10217 24452 10273 24454
rect 10297 24452 10353 24454
rect 10377 24452 10433 24454
rect 10457 24452 10513 24454
rect 10217 23418 10273 23420
rect 10297 23418 10353 23420
rect 10377 23418 10433 23420
rect 10457 23418 10513 23420
rect 10217 23366 10243 23418
rect 10243 23366 10273 23418
rect 10297 23366 10307 23418
rect 10307 23366 10353 23418
rect 10377 23366 10423 23418
rect 10423 23366 10433 23418
rect 10457 23366 10487 23418
rect 10487 23366 10513 23418
rect 10217 23364 10273 23366
rect 10297 23364 10353 23366
rect 10377 23364 10433 23366
rect 10457 23364 10513 23366
rect 10217 22330 10273 22332
rect 10297 22330 10353 22332
rect 10377 22330 10433 22332
rect 10457 22330 10513 22332
rect 10217 22278 10243 22330
rect 10243 22278 10273 22330
rect 10297 22278 10307 22330
rect 10307 22278 10353 22330
rect 10377 22278 10423 22330
rect 10423 22278 10433 22330
rect 10457 22278 10487 22330
rect 10487 22278 10513 22330
rect 10217 22276 10273 22278
rect 10297 22276 10353 22278
rect 10377 22276 10433 22278
rect 10457 22276 10513 22278
rect 10217 21242 10273 21244
rect 10297 21242 10353 21244
rect 10377 21242 10433 21244
rect 10457 21242 10513 21244
rect 10217 21190 10243 21242
rect 10243 21190 10273 21242
rect 10297 21190 10307 21242
rect 10307 21190 10353 21242
rect 10377 21190 10423 21242
rect 10423 21190 10433 21242
rect 10457 21190 10487 21242
rect 10487 21190 10513 21242
rect 10217 21188 10273 21190
rect 10297 21188 10353 21190
rect 10377 21188 10433 21190
rect 10457 21188 10513 21190
rect 10217 20154 10273 20156
rect 10297 20154 10353 20156
rect 10377 20154 10433 20156
rect 10457 20154 10513 20156
rect 10217 20102 10243 20154
rect 10243 20102 10273 20154
rect 10297 20102 10307 20154
rect 10307 20102 10353 20154
rect 10377 20102 10423 20154
rect 10423 20102 10433 20154
rect 10457 20102 10487 20154
rect 10487 20102 10513 20154
rect 10217 20100 10273 20102
rect 10297 20100 10353 20102
rect 10377 20100 10433 20102
rect 10457 20100 10513 20102
rect 10217 19066 10273 19068
rect 10297 19066 10353 19068
rect 10377 19066 10433 19068
rect 10457 19066 10513 19068
rect 10217 19014 10243 19066
rect 10243 19014 10273 19066
rect 10297 19014 10307 19066
rect 10307 19014 10353 19066
rect 10377 19014 10423 19066
rect 10423 19014 10433 19066
rect 10457 19014 10487 19066
rect 10487 19014 10513 19066
rect 10217 19012 10273 19014
rect 10297 19012 10353 19014
rect 10377 19012 10433 19014
rect 10457 19012 10513 19014
rect 10217 17978 10273 17980
rect 10297 17978 10353 17980
rect 10377 17978 10433 17980
rect 10457 17978 10513 17980
rect 10217 17926 10243 17978
rect 10243 17926 10273 17978
rect 10297 17926 10307 17978
rect 10307 17926 10353 17978
rect 10377 17926 10423 17978
rect 10423 17926 10433 17978
rect 10457 17926 10487 17978
rect 10487 17926 10513 17978
rect 10217 17924 10273 17926
rect 10297 17924 10353 17926
rect 10377 17924 10433 17926
rect 10457 17924 10513 17926
rect 10217 16890 10273 16892
rect 10297 16890 10353 16892
rect 10377 16890 10433 16892
rect 10457 16890 10513 16892
rect 10217 16838 10243 16890
rect 10243 16838 10273 16890
rect 10297 16838 10307 16890
rect 10307 16838 10353 16890
rect 10377 16838 10423 16890
rect 10423 16838 10433 16890
rect 10457 16838 10487 16890
rect 10487 16838 10513 16890
rect 10217 16836 10273 16838
rect 10297 16836 10353 16838
rect 10377 16836 10433 16838
rect 10457 16836 10513 16838
rect 10217 15802 10273 15804
rect 10297 15802 10353 15804
rect 10377 15802 10433 15804
rect 10457 15802 10513 15804
rect 10217 15750 10243 15802
rect 10243 15750 10273 15802
rect 10297 15750 10307 15802
rect 10307 15750 10353 15802
rect 10377 15750 10423 15802
rect 10423 15750 10433 15802
rect 10457 15750 10487 15802
rect 10487 15750 10513 15802
rect 10217 15748 10273 15750
rect 10297 15748 10353 15750
rect 10377 15748 10433 15750
rect 10457 15748 10513 15750
rect 14848 29402 14904 29404
rect 14928 29402 14984 29404
rect 15008 29402 15064 29404
rect 15088 29402 15144 29404
rect 14848 29350 14874 29402
rect 14874 29350 14904 29402
rect 14928 29350 14938 29402
rect 14938 29350 14984 29402
rect 15008 29350 15054 29402
rect 15054 29350 15064 29402
rect 15088 29350 15118 29402
rect 15118 29350 15144 29402
rect 14848 29348 14904 29350
rect 14928 29348 14984 29350
rect 15008 29348 15064 29350
rect 15088 29348 15144 29350
rect 24109 29402 24165 29404
rect 24189 29402 24245 29404
rect 24269 29402 24325 29404
rect 24349 29402 24405 29404
rect 24109 29350 24135 29402
rect 24135 29350 24165 29402
rect 24189 29350 24199 29402
rect 24199 29350 24245 29402
rect 24269 29350 24315 29402
rect 24315 29350 24325 29402
rect 24349 29350 24379 29402
rect 24379 29350 24405 29402
rect 24109 29348 24165 29350
rect 24189 29348 24245 29350
rect 24269 29348 24325 29350
rect 24349 29348 24405 29350
rect 19478 28858 19534 28860
rect 19558 28858 19614 28860
rect 19638 28858 19694 28860
rect 19718 28858 19774 28860
rect 19478 28806 19504 28858
rect 19504 28806 19534 28858
rect 19558 28806 19568 28858
rect 19568 28806 19614 28858
rect 19638 28806 19684 28858
rect 19684 28806 19694 28858
rect 19718 28806 19748 28858
rect 19748 28806 19774 28858
rect 19478 28804 19534 28806
rect 19558 28804 19614 28806
rect 19638 28804 19694 28806
rect 19718 28804 19774 28806
rect 14848 28314 14904 28316
rect 14928 28314 14984 28316
rect 15008 28314 15064 28316
rect 15088 28314 15144 28316
rect 14848 28262 14874 28314
rect 14874 28262 14904 28314
rect 14928 28262 14938 28314
rect 14938 28262 14984 28314
rect 15008 28262 15054 28314
rect 15054 28262 15064 28314
rect 15088 28262 15118 28314
rect 15118 28262 15144 28314
rect 14848 28260 14904 28262
rect 14928 28260 14984 28262
rect 15008 28260 15064 28262
rect 15088 28260 15144 28262
rect 24109 28314 24165 28316
rect 24189 28314 24245 28316
rect 24269 28314 24325 28316
rect 24349 28314 24405 28316
rect 24109 28262 24135 28314
rect 24135 28262 24165 28314
rect 24189 28262 24199 28314
rect 24199 28262 24245 28314
rect 24269 28262 24315 28314
rect 24315 28262 24325 28314
rect 24349 28262 24379 28314
rect 24379 28262 24405 28314
rect 24109 28260 24165 28262
rect 24189 28260 24245 28262
rect 24269 28260 24325 28262
rect 24349 28260 24405 28262
rect 19478 27770 19534 27772
rect 19558 27770 19614 27772
rect 19638 27770 19694 27772
rect 19718 27770 19774 27772
rect 19478 27718 19504 27770
rect 19504 27718 19534 27770
rect 19558 27718 19568 27770
rect 19568 27718 19614 27770
rect 19638 27718 19684 27770
rect 19684 27718 19694 27770
rect 19718 27718 19748 27770
rect 19748 27718 19774 27770
rect 19478 27716 19534 27718
rect 19558 27716 19614 27718
rect 19638 27716 19694 27718
rect 19718 27716 19774 27718
rect 14848 27226 14904 27228
rect 14928 27226 14984 27228
rect 15008 27226 15064 27228
rect 15088 27226 15144 27228
rect 14848 27174 14874 27226
rect 14874 27174 14904 27226
rect 14928 27174 14938 27226
rect 14938 27174 14984 27226
rect 15008 27174 15054 27226
rect 15054 27174 15064 27226
rect 15088 27174 15118 27226
rect 15118 27174 15144 27226
rect 14848 27172 14904 27174
rect 14928 27172 14984 27174
rect 15008 27172 15064 27174
rect 15088 27172 15144 27174
rect 24109 27226 24165 27228
rect 24189 27226 24245 27228
rect 24269 27226 24325 27228
rect 24349 27226 24405 27228
rect 24109 27174 24135 27226
rect 24135 27174 24165 27226
rect 24189 27174 24199 27226
rect 24199 27174 24245 27226
rect 24269 27174 24315 27226
rect 24315 27174 24325 27226
rect 24349 27174 24379 27226
rect 24379 27174 24405 27226
rect 24109 27172 24165 27174
rect 24189 27172 24245 27174
rect 24269 27172 24325 27174
rect 24349 27172 24405 27174
rect 19478 26682 19534 26684
rect 19558 26682 19614 26684
rect 19638 26682 19694 26684
rect 19718 26682 19774 26684
rect 19478 26630 19504 26682
rect 19504 26630 19534 26682
rect 19558 26630 19568 26682
rect 19568 26630 19614 26682
rect 19638 26630 19684 26682
rect 19684 26630 19694 26682
rect 19718 26630 19748 26682
rect 19748 26630 19774 26682
rect 19478 26628 19534 26630
rect 19558 26628 19614 26630
rect 19638 26628 19694 26630
rect 19718 26628 19774 26630
rect 14848 26138 14904 26140
rect 14928 26138 14984 26140
rect 15008 26138 15064 26140
rect 15088 26138 15144 26140
rect 14848 26086 14874 26138
rect 14874 26086 14904 26138
rect 14928 26086 14938 26138
rect 14938 26086 14984 26138
rect 15008 26086 15054 26138
rect 15054 26086 15064 26138
rect 15088 26086 15118 26138
rect 15118 26086 15144 26138
rect 14848 26084 14904 26086
rect 14928 26084 14984 26086
rect 15008 26084 15064 26086
rect 15088 26084 15144 26086
rect 24109 26138 24165 26140
rect 24189 26138 24245 26140
rect 24269 26138 24325 26140
rect 24349 26138 24405 26140
rect 24109 26086 24135 26138
rect 24135 26086 24165 26138
rect 24189 26086 24199 26138
rect 24199 26086 24245 26138
rect 24269 26086 24315 26138
rect 24315 26086 24325 26138
rect 24349 26086 24379 26138
rect 24379 26086 24405 26138
rect 24109 26084 24165 26086
rect 24189 26084 24245 26086
rect 24269 26084 24325 26086
rect 24349 26084 24405 26086
rect 19478 25594 19534 25596
rect 19558 25594 19614 25596
rect 19638 25594 19694 25596
rect 19718 25594 19774 25596
rect 19478 25542 19504 25594
rect 19504 25542 19534 25594
rect 19558 25542 19568 25594
rect 19568 25542 19614 25594
rect 19638 25542 19684 25594
rect 19684 25542 19694 25594
rect 19718 25542 19748 25594
rect 19748 25542 19774 25594
rect 19478 25540 19534 25542
rect 19558 25540 19614 25542
rect 19638 25540 19694 25542
rect 19718 25540 19774 25542
rect 14848 25050 14904 25052
rect 14928 25050 14984 25052
rect 15008 25050 15064 25052
rect 15088 25050 15144 25052
rect 14848 24998 14874 25050
rect 14874 24998 14904 25050
rect 14928 24998 14938 25050
rect 14938 24998 14984 25050
rect 15008 24998 15054 25050
rect 15054 24998 15064 25050
rect 15088 24998 15118 25050
rect 15118 24998 15144 25050
rect 14848 24996 14904 24998
rect 14928 24996 14984 24998
rect 15008 24996 15064 24998
rect 15088 24996 15144 24998
rect 24109 25050 24165 25052
rect 24189 25050 24245 25052
rect 24269 25050 24325 25052
rect 24349 25050 24405 25052
rect 24109 24998 24135 25050
rect 24135 24998 24165 25050
rect 24189 24998 24199 25050
rect 24199 24998 24245 25050
rect 24269 24998 24315 25050
rect 24315 24998 24325 25050
rect 24349 24998 24379 25050
rect 24379 24998 24405 25050
rect 24109 24996 24165 24998
rect 24189 24996 24245 24998
rect 24269 24996 24325 24998
rect 24349 24996 24405 24998
rect 19478 24506 19534 24508
rect 19558 24506 19614 24508
rect 19638 24506 19694 24508
rect 19718 24506 19774 24508
rect 19478 24454 19504 24506
rect 19504 24454 19534 24506
rect 19558 24454 19568 24506
rect 19568 24454 19614 24506
rect 19638 24454 19684 24506
rect 19684 24454 19694 24506
rect 19718 24454 19748 24506
rect 19748 24454 19774 24506
rect 19478 24452 19534 24454
rect 19558 24452 19614 24454
rect 19638 24452 19694 24454
rect 19718 24452 19774 24454
rect 14848 23962 14904 23964
rect 14928 23962 14984 23964
rect 15008 23962 15064 23964
rect 15088 23962 15144 23964
rect 14848 23910 14874 23962
rect 14874 23910 14904 23962
rect 14928 23910 14938 23962
rect 14938 23910 14984 23962
rect 15008 23910 15054 23962
rect 15054 23910 15064 23962
rect 15088 23910 15118 23962
rect 15118 23910 15144 23962
rect 14848 23908 14904 23910
rect 14928 23908 14984 23910
rect 15008 23908 15064 23910
rect 15088 23908 15144 23910
rect 24109 23962 24165 23964
rect 24189 23962 24245 23964
rect 24269 23962 24325 23964
rect 24349 23962 24405 23964
rect 24109 23910 24135 23962
rect 24135 23910 24165 23962
rect 24189 23910 24199 23962
rect 24199 23910 24245 23962
rect 24269 23910 24315 23962
rect 24315 23910 24325 23962
rect 24349 23910 24379 23962
rect 24379 23910 24405 23962
rect 24109 23908 24165 23910
rect 24189 23908 24245 23910
rect 24269 23908 24325 23910
rect 24349 23908 24405 23910
rect 19478 23418 19534 23420
rect 19558 23418 19614 23420
rect 19638 23418 19694 23420
rect 19718 23418 19774 23420
rect 19478 23366 19504 23418
rect 19504 23366 19534 23418
rect 19558 23366 19568 23418
rect 19568 23366 19614 23418
rect 19638 23366 19684 23418
rect 19684 23366 19694 23418
rect 19718 23366 19748 23418
rect 19748 23366 19774 23418
rect 19478 23364 19534 23366
rect 19558 23364 19614 23366
rect 19638 23364 19694 23366
rect 19718 23364 19774 23366
rect 14848 22874 14904 22876
rect 14928 22874 14984 22876
rect 15008 22874 15064 22876
rect 15088 22874 15144 22876
rect 14848 22822 14874 22874
rect 14874 22822 14904 22874
rect 14928 22822 14938 22874
rect 14938 22822 14984 22874
rect 15008 22822 15054 22874
rect 15054 22822 15064 22874
rect 15088 22822 15118 22874
rect 15118 22822 15144 22874
rect 14848 22820 14904 22822
rect 14928 22820 14984 22822
rect 15008 22820 15064 22822
rect 15088 22820 15144 22822
rect 24109 22874 24165 22876
rect 24189 22874 24245 22876
rect 24269 22874 24325 22876
rect 24349 22874 24405 22876
rect 24109 22822 24135 22874
rect 24135 22822 24165 22874
rect 24189 22822 24199 22874
rect 24199 22822 24245 22874
rect 24269 22822 24315 22874
rect 24315 22822 24325 22874
rect 24349 22822 24379 22874
rect 24379 22822 24405 22874
rect 24109 22820 24165 22822
rect 24189 22820 24245 22822
rect 24269 22820 24325 22822
rect 24349 22820 24405 22822
rect 19478 22330 19534 22332
rect 19558 22330 19614 22332
rect 19638 22330 19694 22332
rect 19718 22330 19774 22332
rect 19478 22278 19504 22330
rect 19504 22278 19534 22330
rect 19558 22278 19568 22330
rect 19568 22278 19614 22330
rect 19638 22278 19684 22330
rect 19684 22278 19694 22330
rect 19718 22278 19748 22330
rect 19748 22278 19774 22330
rect 19478 22276 19534 22278
rect 19558 22276 19614 22278
rect 19638 22276 19694 22278
rect 19718 22276 19774 22278
rect 14848 21786 14904 21788
rect 14928 21786 14984 21788
rect 15008 21786 15064 21788
rect 15088 21786 15144 21788
rect 14848 21734 14874 21786
rect 14874 21734 14904 21786
rect 14928 21734 14938 21786
rect 14938 21734 14984 21786
rect 15008 21734 15054 21786
rect 15054 21734 15064 21786
rect 15088 21734 15118 21786
rect 15118 21734 15144 21786
rect 14848 21732 14904 21734
rect 14928 21732 14984 21734
rect 15008 21732 15064 21734
rect 15088 21732 15144 21734
rect 24109 21786 24165 21788
rect 24189 21786 24245 21788
rect 24269 21786 24325 21788
rect 24349 21786 24405 21788
rect 24109 21734 24135 21786
rect 24135 21734 24165 21786
rect 24189 21734 24199 21786
rect 24199 21734 24245 21786
rect 24269 21734 24315 21786
rect 24315 21734 24325 21786
rect 24349 21734 24379 21786
rect 24379 21734 24405 21786
rect 24109 21732 24165 21734
rect 24189 21732 24245 21734
rect 24269 21732 24325 21734
rect 24349 21732 24405 21734
rect 19478 21242 19534 21244
rect 19558 21242 19614 21244
rect 19638 21242 19694 21244
rect 19718 21242 19774 21244
rect 19478 21190 19504 21242
rect 19504 21190 19534 21242
rect 19558 21190 19568 21242
rect 19568 21190 19614 21242
rect 19638 21190 19684 21242
rect 19684 21190 19694 21242
rect 19718 21190 19748 21242
rect 19748 21190 19774 21242
rect 19478 21188 19534 21190
rect 19558 21188 19614 21190
rect 19638 21188 19694 21190
rect 19718 21188 19774 21190
rect 14848 20698 14904 20700
rect 14928 20698 14984 20700
rect 15008 20698 15064 20700
rect 15088 20698 15144 20700
rect 14848 20646 14874 20698
rect 14874 20646 14904 20698
rect 14928 20646 14938 20698
rect 14938 20646 14984 20698
rect 15008 20646 15054 20698
rect 15054 20646 15064 20698
rect 15088 20646 15118 20698
rect 15118 20646 15144 20698
rect 14848 20644 14904 20646
rect 14928 20644 14984 20646
rect 15008 20644 15064 20646
rect 15088 20644 15144 20646
rect 24109 20698 24165 20700
rect 24189 20698 24245 20700
rect 24269 20698 24325 20700
rect 24349 20698 24405 20700
rect 24109 20646 24135 20698
rect 24135 20646 24165 20698
rect 24189 20646 24199 20698
rect 24199 20646 24245 20698
rect 24269 20646 24315 20698
rect 24315 20646 24325 20698
rect 24349 20646 24379 20698
rect 24379 20646 24405 20698
rect 24109 20644 24165 20646
rect 24189 20644 24245 20646
rect 24269 20644 24325 20646
rect 24349 20644 24405 20646
rect 19478 20154 19534 20156
rect 19558 20154 19614 20156
rect 19638 20154 19694 20156
rect 19718 20154 19774 20156
rect 19478 20102 19504 20154
rect 19504 20102 19534 20154
rect 19558 20102 19568 20154
rect 19568 20102 19614 20154
rect 19638 20102 19684 20154
rect 19684 20102 19694 20154
rect 19718 20102 19748 20154
rect 19748 20102 19774 20154
rect 19478 20100 19534 20102
rect 19558 20100 19614 20102
rect 19638 20100 19694 20102
rect 19718 20100 19774 20102
rect 14848 19610 14904 19612
rect 14928 19610 14984 19612
rect 15008 19610 15064 19612
rect 15088 19610 15144 19612
rect 14848 19558 14874 19610
rect 14874 19558 14904 19610
rect 14928 19558 14938 19610
rect 14938 19558 14984 19610
rect 15008 19558 15054 19610
rect 15054 19558 15064 19610
rect 15088 19558 15118 19610
rect 15118 19558 15144 19610
rect 14848 19556 14904 19558
rect 14928 19556 14984 19558
rect 15008 19556 15064 19558
rect 15088 19556 15144 19558
rect 24109 19610 24165 19612
rect 24189 19610 24245 19612
rect 24269 19610 24325 19612
rect 24349 19610 24405 19612
rect 24109 19558 24135 19610
rect 24135 19558 24165 19610
rect 24189 19558 24199 19610
rect 24199 19558 24245 19610
rect 24269 19558 24315 19610
rect 24315 19558 24325 19610
rect 24349 19558 24379 19610
rect 24379 19558 24405 19610
rect 24109 19556 24165 19558
rect 24189 19556 24245 19558
rect 24269 19556 24325 19558
rect 24349 19556 24405 19558
rect 19478 19066 19534 19068
rect 19558 19066 19614 19068
rect 19638 19066 19694 19068
rect 19718 19066 19774 19068
rect 19478 19014 19504 19066
rect 19504 19014 19534 19066
rect 19558 19014 19568 19066
rect 19568 19014 19614 19066
rect 19638 19014 19684 19066
rect 19684 19014 19694 19066
rect 19718 19014 19748 19066
rect 19748 19014 19774 19066
rect 19478 19012 19534 19014
rect 19558 19012 19614 19014
rect 19638 19012 19694 19014
rect 19718 19012 19774 19014
rect 14848 18522 14904 18524
rect 14928 18522 14984 18524
rect 15008 18522 15064 18524
rect 15088 18522 15144 18524
rect 14848 18470 14874 18522
rect 14874 18470 14904 18522
rect 14928 18470 14938 18522
rect 14938 18470 14984 18522
rect 15008 18470 15054 18522
rect 15054 18470 15064 18522
rect 15088 18470 15118 18522
rect 15118 18470 15144 18522
rect 14848 18468 14904 18470
rect 14928 18468 14984 18470
rect 15008 18468 15064 18470
rect 15088 18468 15144 18470
rect 24109 18522 24165 18524
rect 24189 18522 24245 18524
rect 24269 18522 24325 18524
rect 24349 18522 24405 18524
rect 24109 18470 24135 18522
rect 24135 18470 24165 18522
rect 24189 18470 24199 18522
rect 24199 18470 24245 18522
rect 24269 18470 24315 18522
rect 24315 18470 24325 18522
rect 24349 18470 24379 18522
rect 24379 18470 24405 18522
rect 24109 18468 24165 18470
rect 24189 18468 24245 18470
rect 24269 18468 24325 18470
rect 24349 18468 24405 18470
rect 19478 17978 19534 17980
rect 19558 17978 19614 17980
rect 19638 17978 19694 17980
rect 19718 17978 19774 17980
rect 19478 17926 19504 17978
rect 19504 17926 19534 17978
rect 19558 17926 19568 17978
rect 19568 17926 19614 17978
rect 19638 17926 19684 17978
rect 19684 17926 19694 17978
rect 19718 17926 19748 17978
rect 19748 17926 19774 17978
rect 19478 17924 19534 17926
rect 19558 17924 19614 17926
rect 19638 17924 19694 17926
rect 19718 17924 19774 17926
rect 14848 17434 14904 17436
rect 14928 17434 14984 17436
rect 15008 17434 15064 17436
rect 15088 17434 15144 17436
rect 14848 17382 14874 17434
rect 14874 17382 14904 17434
rect 14928 17382 14938 17434
rect 14938 17382 14984 17434
rect 15008 17382 15054 17434
rect 15054 17382 15064 17434
rect 15088 17382 15118 17434
rect 15118 17382 15144 17434
rect 14848 17380 14904 17382
rect 14928 17380 14984 17382
rect 15008 17380 15064 17382
rect 15088 17380 15144 17382
rect 24109 17434 24165 17436
rect 24189 17434 24245 17436
rect 24269 17434 24325 17436
rect 24349 17434 24405 17436
rect 24109 17382 24135 17434
rect 24135 17382 24165 17434
rect 24189 17382 24199 17434
rect 24199 17382 24245 17434
rect 24269 17382 24315 17434
rect 24315 17382 24325 17434
rect 24349 17382 24379 17434
rect 24379 17382 24405 17434
rect 24109 17380 24165 17382
rect 24189 17380 24245 17382
rect 24269 17380 24325 17382
rect 24349 17380 24405 17382
rect 28170 17060 28226 17096
rect 28170 17040 28172 17060
rect 28172 17040 28224 17060
rect 28224 17040 28226 17060
rect 19478 16890 19534 16892
rect 19558 16890 19614 16892
rect 19638 16890 19694 16892
rect 19718 16890 19774 16892
rect 19478 16838 19504 16890
rect 19504 16838 19534 16890
rect 19558 16838 19568 16890
rect 19568 16838 19614 16890
rect 19638 16838 19684 16890
rect 19684 16838 19694 16890
rect 19718 16838 19748 16890
rect 19748 16838 19774 16890
rect 19478 16836 19534 16838
rect 19558 16836 19614 16838
rect 19638 16836 19694 16838
rect 19718 16836 19774 16838
rect 14848 16346 14904 16348
rect 14928 16346 14984 16348
rect 15008 16346 15064 16348
rect 15088 16346 15144 16348
rect 14848 16294 14874 16346
rect 14874 16294 14904 16346
rect 14928 16294 14938 16346
rect 14938 16294 14984 16346
rect 15008 16294 15054 16346
rect 15054 16294 15064 16346
rect 15088 16294 15118 16346
rect 15118 16294 15144 16346
rect 14848 16292 14904 16294
rect 14928 16292 14984 16294
rect 15008 16292 15064 16294
rect 15088 16292 15144 16294
rect 24109 16346 24165 16348
rect 24189 16346 24245 16348
rect 24269 16346 24325 16348
rect 24349 16346 24405 16348
rect 24109 16294 24135 16346
rect 24135 16294 24165 16346
rect 24189 16294 24199 16346
rect 24199 16294 24245 16346
rect 24269 16294 24315 16346
rect 24315 16294 24325 16346
rect 24349 16294 24379 16346
rect 24379 16294 24405 16346
rect 24109 16292 24165 16294
rect 24189 16292 24245 16294
rect 24269 16292 24325 16294
rect 24349 16292 24405 16294
rect 19478 15802 19534 15804
rect 19558 15802 19614 15804
rect 19638 15802 19694 15804
rect 19718 15802 19774 15804
rect 19478 15750 19504 15802
rect 19504 15750 19534 15802
rect 19558 15750 19568 15802
rect 19568 15750 19614 15802
rect 19638 15750 19684 15802
rect 19684 15750 19694 15802
rect 19718 15750 19748 15802
rect 19748 15750 19774 15802
rect 19478 15748 19534 15750
rect 19558 15748 19614 15750
rect 19638 15748 19694 15750
rect 19718 15748 19774 15750
rect 14848 15258 14904 15260
rect 14928 15258 14984 15260
rect 15008 15258 15064 15260
rect 15088 15258 15144 15260
rect 14848 15206 14874 15258
rect 14874 15206 14904 15258
rect 14928 15206 14938 15258
rect 14938 15206 14984 15258
rect 15008 15206 15054 15258
rect 15054 15206 15064 15258
rect 15088 15206 15118 15258
rect 15118 15206 15144 15258
rect 14848 15204 14904 15206
rect 14928 15204 14984 15206
rect 15008 15204 15064 15206
rect 15088 15204 15144 15206
rect 24109 15258 24165 15260
rect 24189 15258 24245 15260
rect 24269 15258 24325 15260
rect 24349 15258 24405 15260
rect 24109 15206 24135 15258
rect 24135 15206 24165 15258
rect 24189 15206 24199 15258
rect 24199 15206 24245 15258
rect 24269 15206 24315 15258
rect 24315 15206 24325 15258
rect 24349 15206 24379 15258
rect 24379 15206 24405 15258
rect 24109 15204 24165 15206
rect 24189 15204 24245 15206
rect 24269 15204 24325 15206
rect 24349 15204 24405 15206
rect 10217 14714 10273 14716
rect 10297 14714 10353 14716
rect 10377 14714 10433 14716
rect 10457 14714 10513 14716
rect 10217 14662 10243 14714
rect 10243 14662 10273 14714
rect 10297 14662 10307 14714
rect 10307 14662 10353 14714
rect 10377 14662 10423 14714
rect 10423 14662 10433 14714
rect 10457 14662 10487 14714
rect 10487 14662 10513 14714
rect 10217 14660 10273 14662
rect 10297 14660 10353 14662
rect 10377 14660 10433 14662
rect 10457 14660 10513 14662
rect 10217 13626 10273 13628
rect 10297 13626 10353 13628
rect 10377 13626 10433 13628
rect 10457 13626 10513 13628
rect 10217 13574 10243 13626
rect 10243 13574 10273 13626
rect 10297 13574 10307 13626
rect 10307 13574 10353 13626
rect 10377 13574 10423 13626
rect 10423 13574 10433 13626
rect 10457 13574 10487 13626
rect 10487 13574 10513 13626
rect 10217 13572 10273 13574
rect 10297 13572 10353 13574
rect 10377 13572 10433 13574
rect 10457 13572 10513 13574
rect 5586 13082 5642 13084
rect 5666 13082 5722 13084
rect 5746 13082 5802 13084
rect 5826 13082 5882 13084
rect 5586 13030 5612 13082
rect 5612 13030 5642 13082
rect 5666 13030 5676 13082
rect 5676 13030 5722 13082
rect 5746 13030 5792 13082
rect 5792 13030 5802 13082
rect 5826 13030 5856 13082
rect 5856 13030 5882 13082
rect 5586 13028 5642 13030
rect 5666 13028 5722 13030
rect 5746 13028 5802 13030
rect 5826 13028 5882 13030
rect 5586 11994 5642 11996
rect 5666 11994 5722 11996
rect 5746 11994 5802 11996
rect 5826 11994 5882 11996
rect 5586 11942 5612 11994
rect 5612 11942 5642 11994
rect 5666 11942 5676 11994
rect 5676 11942 5722 11994
rect 5746 11942 5792 11994
rect 5792 11942 5802 11994
rect 5826 11942 5856 11994
rect 5856 11942 5882 11994
rect 5586 11940 5642 11942
rect 5666 11940 5722 11942
rect 5746 11940 5802 11942
rect 5826 11940 5882 11942
rect 5586 10906 5642 10908
rect 5666 10906 5722 10908
rect 5746 10906 5802 10908
rect 5826 10906 5882 10908
rect 5586 10854 5612 10906
rect 5612 10854 5642 10906
rect 5666 10854 5676 10906
rect 5676 10854 5722 10906
rect 5746 10854 5792 10906
rect 5792 10854 5802 10906
rect 5826 10854 5856 10906
rect 5856 10854 5882 10906
rect 5586 10852 5642 10854
rect 5666 10852 5722 10854
rect 5746 10852 5802 10854
rect 5826 10852 5882 10854
rect 10217 12538 10273 12540
rect 10297 12538 10353 12540
rect 10377 12538 10433 12540
rect 10457 12538 10513 12540
rect 10217 12486 10243 12538
rect 10243 12486 10273 12538
rect 10297 12486 10307 12538
rect 10307 12486 10353 12538
rect 10377 12486 10423 12538
rect 10423 12486 10433 12538
rect 10457 12486 10487 12538
rect 10487 12486 10513 12538
rect 10217 12484 10273 12486
rect 10297 12484 10353 12486
rect 10377 12484 10433 12486
rect 10457 12484 10513 12486
rect 10217 11450 10273 11452
rect 10297 11450 10353 11452
rect 10377 11450 10433 11452
rect 10457 11450 10513 11452
rect 10217 11398 10243 11450
rect 10243 11398 10273 11450
rect 10297 11398 10307 11450
rect 10307 11398 10353 11450
rect 10377 11398 10423 11450
rect 10423 11398 10433 11450
rect 10457 11398 10487 11450
rect 10487 11398 10513 11450
rect 10217 11396 10273 11398
rect 10297 11396 10353 11398
rect 10377 11396 10433 11398
rect 10457 11396 10513 11398
rect 10217 10362 10273 10364
rect 10297 10362 10353 10364
rect 10377 10362 10433 10364
rect 10457 10362 10513 10364
rect 10217 10310 10243 10362
rect 10243 10310 10273 10362
rect 10297 10310 10307 10362
rect 10307 10310 10353 10362
rect 10377 10310 10423 10362
rect 10423 10310 10433 10362
rect 10457 10310 10487 10362
rect 10487 10310 10513 10362
rect 10217 10308 10273 10310
rect 10297 10308 10353 10310
rect 10377 10308 10433 10310
rect 10457 10308 10513 10310
rect 5586 9818 5642 9820
rect 5666 9818 5722 9820
rect 5746 9818 5802 9820
rect 5826 9818 5882 9820
rect 5586 9766 5612 9818
rect 5612 9766 5642 9818
rect 5666 9766 5676 9818
rect 5676 9766 5722 9818
rect 5746 9766 5792 9818
rect 5792 9766 5802 9818
rect 5826 9766 5856 9818
rect 5856 9766 5882 9818
rect 5586 9764 5642 9766
rect 5666 9764 5722 9766
rect 5746 9764 5802 9766
rect 5826 9764 5882 9766
rect 10217 9274 10273 9276
rect 10297 9274 10353 9276
rect 10377 9274 10433 9276
rect 10457 9274 10513 9276
rect 10217 9222 10243 9274
rect 10243 9222 10273 9274
rect 10297 9222 10307 9274
rect 10307 9222 10353 9274
rect 10377 9222 10423 9274
rect 10423 9222 10433 9274
rect 10457 9222 10487 9274
rect 10487 9222 10513 9274
rect 10217 9220 10273 9222
rect 10297 9220 10353 9222
rect 10377 9220 10433 9222
rect 10457 9220 10513 9222
rect 5586 8730 5642 8732
rect 5666 8730 5722 8732
rect 5746 8730 5802 8732
rect 5826 8730 5882 8732
rect 5586 8678 5612 8730
rect 5612 8678 5642 8730
rect 5666 8678 5676 8730
rect 5676 8678 5722 8730
rect 5746 8678 5792 8730
rect 5792 8678 5802 8730
rect 5826 8678 5856 8730
rect 5856 8678 5882 8730
rect 5586 8676 5642 8678
rect 5666 8676 5722 8678
rect 5746 8676 5802 8678
rect 5826 8676 5882 8678
rect 5586 7642 5642 7644
rect 5666 7642 5722 7644
rect 5746 7642 5802 7644
rect 5826 7642 5882 7644
rect 5586 7590 5612 7642
rect 5612 7590 5642 7642
rect 5666 7590 5676 7642
rect 5676 7590 5722 7642
rect 5746 7590 5792 7642
rect 5792 7590 5802 7642
rect 5826 7590 5856 7642
rect 5856 7590 5882 7642
rect 5586 7588 5642 7590
rect 5666 7588 5722 7590
rect 5746 7588 5802 7590
rect 5826 7588 5882 7590
rect 5586 6554 5642 6556
rect 5666 6554 5722 6556
rect 5746 6554 5802 6556
rect 5826 6554 5882 6556
rect 5586 6502 5612 6554
rect 5612 6502 5642 6554
rect 5666 6502 5676 6554
rect 5676 6502 5722 6554
rect 5746 6502 5792 6554
rect 5792 6502 5802 6554
rect 5826 6502 5856 6554
rect 5856 6502 5882 6554
rect 5586 6500 5642 6502
rect 5666 6500 5722 6502
rect 5746 6500 5802 6502
rect 5826 6500 5882 6502
rect 10217 8186 10273 8188
rect 10297 8186 10353 8188
rect 10377 8186 10433 8188
rect 10457 8186 10513 8188
rect 10217 8134 10243 8186
rect 10243 8134 10273 8186
rect 10297 8134 10307 8186
rect 10307 8134 10353 8186
rect 10377 8134 10423 8186
rect 10423 8134 10433 8186
rect 10457 8134 10487 8186
rect 10487 8134 10513 8186
rect 10217 8132 10273 8134
rect 10297 8132 10353 8134
rect 10377 8132 10433 8134
rect 10457 8132 10513 8134
rect 10217 7098 10273 7100
rect 10297 7098 10353 7100
rect 10377 7098 10433 7100
rect 10457 7098 10513 7100
rect 10217 7046 10243 7098
rect 10243 7046 10273 7098
rect 10297 7046 10307 7098
rect 10307 7046 10353 7098
rect 10377 7046 10423 7098
rect 10423 7046 10433 7098
rect 10457 7046 10487 7098
rect 10487 7046 10513 7098
rect 10217 7044 10273 7046
rect 10297 7044 10353 7046
rect 10377 7044 10433 7046
rect 10457 7044 10513 7046
rect 10217 6010 10273 6012
rect 10297 6010 10353 6012
rect 10377 6010 10433 6012
rect 10457 6010 10513 6012
rect 10217 5958 10243 6010
rect 10243 5958 10273 6010
rect 10297 5958 10307 6010
rect 10307 5958 10353 6010
rect 10377 5958 10423 6010
rect 10423 5958 10433 6010
rect 10457 5958 10487 6010
rect 10487 5958 10513 6010
rect 10217 5956 10273 5958
rect 10297 5956 10353 5958
rect 10377 5956 10433 5958
rect 10457 5956 10513 5958
rect 5586 5466 5642 5468
rect 5666 5466 5722 5468
rect 5746 5466 5802 5468
rect 5826 5466 5882 5468
rect 5586 5414 5612 5466
rect 5612 5414 5642 5466
rect 5666 5414 5676 5466
rect 5676 5414 5722 5466
rect 5746 5414 5792 5466
rect 5792 5414 5802 5466
rect 5826 5414 5856 5466
rect 5856 5414 5882 5466
rect 5586 5412 5642 5414
rect 5666 5412 5722 5414
rect 5746 5412 5802 5414
rect 5826 5412 5882 5414
rect 10217 4922 10273 4924
rect 10297 4922 10353 4924
rect 10377 4922 10433 4924
rect 10457 4922 10513 4924
rect 10217 4870 10243 4922
rect 10243 4870 10273 4922
rect 10297 4870 10307 4922
rect 10307 4870 10353 4922
rect 10377 4870 10423 4922
rect 10423 4870 10433 4922
rect 10457 4870 10487 4922
rect 10487 4870 10513 4922
rect 10217 4868 10273 4870
rect 10297 4868 10353 4870
rect 10377 4868 10433 4870
rect 10457 4868 10513 4870
rect 5586 4378 5642 4380
rect 5666 4378 5722 4380
rect 5746 4378 5802 4380
rect 5826 4378 5882 4380
rect 5586 4326 5612 4378
rect 5612 4326 5642 4378
rect 5666 4326 5676 4378
rect 5676 4326 5722 4378
rect 5746 4326 5792 4378
rect 5792 4326 5802 4378
rect 5826 4326 5856 4378
rect 5856 4326 5882 4378
rect 5586 4324 5642 4326
rect 5666 4324 5722 4326
rect 5746 4324 5802 4326
rect 5826 4324 5882 4326
rect 10217 3834 10273 3836
rect 10297 3834 10353 3836
rect 10377 3834 10433 3836
rect 10457 3834 10513 3836
rect 10217 3782 10243 3834
rect 10243 3782 10273 3834
rect 10297 3782 10307 3834
rect 10307 3782 10353 3834
rect 10377 3782 10423 3834
rect 10423 3782 10433 3834
rect 10457 3782 10487 3834
rect 10487 3782 10513 3834
rect 10217 3780 10273 3782
rect 10297 3780 10353 3782
rect 10377 3780 10433 3782
rect 10457 3780 10513 3782
rect 5586 3290 5642 3292
rect 5666 3290 5722 3292
rect 5746 3290 5802 3292
rect 5826 3290 5882 3292
rect 5586 3238 5612 3290
rect 5612 3238 5642 3290
rect 5666 3238 5676 3290
rect 5676 3238 5722 3290
rect 5746 3238 5792 3290
rect 5792 3238 5802 3290
rect 5826 3238 5856 3290
rect 5856 3238 5882 3290
rect 5586 3236 5642 3238
rect 5666 3236 5722 3238
rect 5746 3236 5802 3238
rect 5826 3236 5882 3238
rect 10217 2746 10273 2748
rect 10297 2746 10353 2748
rect 10377 2746 10433 2748
rect 10457 2746 10513 2748
rect 10217 2694 10243 2746
rect 10243 2694 10273 2746
rect 10297 2694 10307 2746
rect 10307 2694 10353 2746
rect 10377 2694 10423 2746
rect 10423 2694 10433 2746
rect 10457 2694 10487 2746
rect 10487 2694 10513 2746
rect 10217 2692 10273 2694
rect 10297 2692 10353 2694
rect 10377 2692 10433 2694
rect 10457 2692 10513 2694
rect 5586 2202 5642 2204
rect 5666 2202 5722 2204
rect 5746 2202 5802 2204
rect 5826 2202 5882 2204
rect 5586 2150 5612 2202
rect 5612 2150 5642 2202
rect 5666 2150 5676 2202
rect 5676 2150 5722 2202
rect 5746 2150 5792 2202
rect 5792 2150 5802 2202
rect 5826 2150 5856 2202
rect 5856 2150 5882 2202
rect 5586 2148 5642 2150
rect 5666 2148 5722 2150
rect 5746 2148 5802 2150
rect 5826 2148 5882 2150
rect 19478 14714 19534 14716
rect 19558 14714 19614 14716
rect 19638 14714 19694 14716
rect 19718 14714 19774 14716
rect 19478 14662 19504 14714
rect 19504 14662 19534 14714
rect 19558 14662 19568 14714
rect 19568 14662 19614 14714
rect 19638 14662 19684 14714
rect 19684 14662 19694 14714
rect 19718 14662 19748 14714
rect 19748 14662 19774 14714
rect 19478 14660 19534 14662
rect 19558 14660 19614 14662
rect 19638 14660 19694 14662
rect 19718 14660 19774 14662
rect 14848 14170 14904 14172
rect 14928 14170 14984 14172
rect 15008 14170 15064 14172
rect 15088 14170 15144 14172
rect 14848 14118 14874 14170
rect 14874 14118 14904 14170
rect 14928 14118 14938 14170
rect 14938 14118 14984 14170
rect 15008 14118 15054 14170
rect 15054 14118 15064 14170
rect 15088 14118 15118 14170
rect 15118 14118 15144 14170
rect 14848 14116 14904 14118
rect 14928 14116 14984 14118
rect 15008 14116 15064 14118
rect 15088 14116 15144 14118
rect 24109 14170 24165 14172
rect 24189 14170 24245 14172
rect 24269 14170 24325 14172
rect 24349 14170 24405 14172
rect 24109 14118 24135 14170
rect 24135 14118 24165 14170
rect 24189 14118 24199 14170
rect 24199 14118 24245 14170
rect 24269 14118 24315 14170
rect 24315 14118 24325 14170
rect 24349 14118 24379 14170
rect 24379 14118 24405 14170
rect 24109 14116 24165 14118
rect 24189 14116 24245 14118
rect 24269 14116 24325 14118
rect 24349 14116 24405 14118
rect 19478 13626 19534 13628
rect 19558 13626 19614 13628
rect 19638 13626 19694 13628
rect 19718 13626 19774 13628
rect 19478 13574 19504 13626
rect 19504 13574 19534 13626
rect 19558 13574 19568 13626
rect 19568 13574 19614 13626
rect 19638 13574 19684 13626
rect 19684 13574 19694 13626
rect 19718 13574 19748 13626
rect 19748 13574 19774 13626
rect 19478 13572 19534 13574
rect 19558 13572 19614 13574
rect 19638 13572 19694 13574
rect 19718 13572 19774 13574
rect 14848 13082 14904 13084
rect 14928 13082 14984 13084
rect 15008 13082 15064 13084
rect 15088 13082 15144 13084
rect 14848 13030 14874 13082
rect 14874 13030 14904 13082
rect 14928 13030 14938 13082
rect 14938 13030 14984 13082
rect 15008 13030 15054 13082
rect 15054 13030 15064 13082
rect 15088 13030 15118 13082
rect 15118 13030 15144 13082
rect 14848 13028 14904 13030
rect 14928 13028 14984 13030
rect 15008 13028 15064 13030
rect 15088 13028 15144 13030
rect 24109 13082 24165 13084
rect 24189 13082 24245 13084
rect 24269 13082 24325 13084
rect 24349 13082 24405 13084
rect 24109 13030 24135 13082
rect 24135 13030 24165 13082
rect 24189 13030 24199 13082
rect 24199 13030 24245 13082
rect 24269 13030 24315 13082
rect 24315 13030 24325 13082
rect 24349 13030 24379 13082
rect 24379 13030 24405 13082
rect 24109 13028 24165 13030
rect 24189 13028 24245 13030
rect 24269 13028 24325 13030
rect 24349 13028 24405 13030
rect 19478 12538 19534 12540
rect 19558 12538 19614 12540
rect 19638 12538 19694 12540
rect 19718 12538 19774 12540
rect 19478 12486 19504 12538
rect 19504 12486 19534 12538
rect 19558 12486 19568 12538
rect 19568 12486 19614 12538
rect 19638 12486 19684 12538
rect 19684 12486 19694 12538
rect 19718 12486 19748 12538
rect 19748 12486 19774 12538
rect 19478 12484 19534 12486
rect 19558 12484 19614 12486
rect 19638 12484 19694 12486
rect 19718 12484 19774 12486
rect 14848 11994 14904 11996
rect 14928 11994 14984 11996
rect 15008 11994 15064 11996
rect 15088 11994 15144 11996
rect 14848 11942 14874 11994
rect 14874 11942 14904 11994
rect 14928 11942 14938 11994
rect 14938 11942 14984 11994
rect 15008 11942 15054 11994
rect 15054 11942 15064 11994
rect 15088 11942 15118 11994
rect 15118 11942 15144 11994
rect 14848 11940 14904 11942
rect 14928 11940 14984 11942
rect 15008 11940 15064 11942
rect 15088 11940 15144 11942
rect 24109 11994 24165 11996
rect 24189 11994 24245 11996
rect 24269 11994 24325 11996
rect 24349 11994 24405 11996
rect 24109 11942 24135 11994
rect 24135 11942 24165 11994
rect 24189 11942 24199 11994
rect 24199 11942 24245 11994
rect 24269 11942 24315 11994
rect 24315 11942 24325 11994
rect 24349 11942 24379 11994
rect 24379 11942 24405 11994
rect 24109 11940 24165 11942
rect 24189 11940 24245 11942
rect 24269 11940 24325 11942
rect 24349 11940 24405 11942
rect 14848 10906 14904 10908
rect 14928 10906 14984 10908
rect 15008 10906 15064 10908
rect 15088 10906 15144 10908
rect 14848 10854 14874 10906
rect 14874 10854 14904 10906
rect 14928 10854 14938 10906
rect 14938 10854 14984 10906
rect 15008 10854 15054 10906
rect 15054 10854 15064 10906
rect 15088 10854 15118 10906
rect 15118 10854 15144 10906
rect 14848 10852 14904 10854
rect 14928 10852 14984 10854
rect 15008 10852 15064 10854
rect 15088 10852 15144 10854
rect 19478 11450 19534 11452
rect 19558 11450 19614 11452
rect 19638 11450 19694 11452
rect 19718 11450 19774 11452
rect 19478 11398 19504 11450
rect 19504 11398 19534 11450
rect 19558 11398 19568 11450
rect 19568 11398 19614 11450
rect 19638 11398 19684 11450
rect 19684 11398 19694 11450
rect 19718 11398 19748 11450
rect 19748 11398 19774 11450
rect 19478 11396 19534 11398
rect 19558 11396 19614 11398
rect 19638 11396 19694 11398
rect 19718 11396 19774 11398
rect 24109 10906 24165 10908
rect 24189 10906 24245 10908
rect 24269 10906 24325 10908
rect 24349 10906 24405 10908
rect 24109 10854 24135 10906
rect 24135 10854 24165 10906
rect 24189 10854 24199 10906
rect 24199 10854 24245 10906
rect 24269 10854 24315 10906
rect 24315 10854 24325 10906
rect 24349 10854 24379 10906
rect 24379 10854 24405 10906
rect 24109 10852 24165 10854
rect 24189 10852 24245 10854
rect 24269 10852 24325 10854
rect 24349 10852 24405 10854
rect 19478 10362 19534 10364
rect 19558 10362 19614 10364
rect 19638 10362 19694 10364
rect 19718 10362 19774 10364
rect 19478 10310 19504 10362
rect 19504 10310 19534 10362
rect 19558 10310 19568 10362
rect 19568 10310 19614 10362
rect 19638 10310 19684 10362
rect 19684 10310 19694 10362
rect 19718 10310 19748 10362
rect 19748 10310 19774 10362
rect 19478 10308 19534 10310
rect 19558 10308 19614 10310
rect 19638 10308 19694 10310
rect 19718 10308 19774 10310
rect 14848 9818 14904 9820
rect 14928 9818 14984 9820
rect 15008 9818 15064 9820
rect 15088 9818 15144 9820
rect 14848 9766 14874 9818
rect 14874 9766 14904 9818
rect 14928 9766 14938 9818
rect 14938 9766 14984 9818
rect 15008 9766 15054 9818
rect 15054 9766 15064 9818
rect 15088 9766 15118 9818
rect 15118 9766 15144 9818
rect 14848 9764 14904 9766
rect 14928 9764 14984 9766
rect 15008 9764 15064 9766
rect 15088 9764 15144 9766
rect 24109 9818 24165 9820
rect 24189 9818 24245 9820
rect 24269 9818 24325 9820
rect 24349 9818 24405 9820
rect 24109 9766 24135 9818
rect 24135 9766 24165 9818
rect 24189 9766 24199 9818
rect 24199 9766 24245 9818
rect 24269 9766 24315 9818
rect 24315 9766 24325 9818
rect 24349 9766 24379 9818
rect 24379 9766 24405 9818
rect 24109 9764 24165 9766
rect 24189 9764 24245 9766
rect 24269 9764 24325 9766
rect 24349 9764 24405 9766
rect 14848 8730 14904 8732
rect 14928 8730 14984 8732
rect 15008 8730 15064 8732
rect 15088 8730 15144 8732
rect 14848 8678 14874 8730
rect 14874 8678 14904 8730
rect 14928 8678 14938 8730
rect 14938 8678 14984 8730
rect 15008 8678 15054 8730
rect 15054 8678 15064 8730
rect 15088 8678 15118 8730
rect 15118 8678 15144 8730
rect 14848 8676 14904 8678
rect 14928 8676 14984 8678
rect 15008 8676 15064 8678
rect 15088 8676 15144 8678
rect 19478 9274 19534 9276
rect 19558 9274 19614 9276
rect 19638 9274 19694 9276
rect 19718 9274 19774 9276
rect 19478 9222 19504 9274
rect 19504 9222 19534 9274
rect 19558 9222 19568 9274
rect 19568 9222 19614 9274
rect 19638 9222 19684 9274
rect 19684 9222 19694 9274
rect 19718 9222 19748 9274
rect 19748 9222 19774 9274
rect 19478 9220 19534 9222
rect 19558 9220 19614 9222
rect 19638 9220 19694 9222
rect 19718 9220 19774 9222
rect 24109 8730 24165 8732
rect 24189 8730 24245 8732
rect 24269 8730 24325 8732
rect 24349 8730 24405 8732
rect 24109 8678 24135 8730
rect 24135 8678 24165 8730
rect 24189 8678 24199 8730
rect 24199 8678 24245 8730
rect 24269 8678 24315 8730
rect 24315 8678 24325 8730
rect 24349 8678 24379 8730
rect 24379 8678 24405 8730
rect 24109 8676 24165 8678
rect 24189 8676 24245 8678
rect 24269 8676 24325 8678
rect 24349 8676 24405 8678
rect 19478 8186 19534 8188
rect 19558 8186 19614 8188
rect 19638 8186 19694 8188
rect 19718 8186 19774 8188
rect 19478 8134 19504 8186
rect 19504 8134 19534 8186
rect 19558 8134 19568 8186
rect 19568 8134 19614 8186
rect 19638 8134 19684 8186
rect 19684 8134 19694 8186
rect 19718 8134 19748 8186
rect 19748 8134 19774 8186
rect 19478 8132 19534 8134
rect 19558 8132 19614 8134
rect 19638 8132 19694 8134
rect 19718 8132 19774 8134
rect 14848 7642 14904 7644
rect 14928 7642 14984 7644
rect 15008 7642 15064 7644
rect 15088 7642 15144 7644
rect 14848 7590 14874 7642
rect 14874 7590 14904 7642
rect 14928 7590 14938 7642
rect 14938 7590 14984 7642
rect 15008 7590 15054 7642
rect 15054 7590 15064 7642
rect 15088 7590 15118 7642
rect 15118 7590 15144 7642
rect 14848 7588 14904 7590
rect 14928 7588 14984 7590
rect 15008 7588 15064 7590
rect 15088 7588 15144 7590
rect 24109 7642 24165 7644
rect 24189 7642 24245 7644
rect 24269 7642 24325 7644
rect 24349 7642 24405 7644
rect 24109 7590 24135 7642
rect 24135 7590 24165 7642
rect 24189 7590 24199 7642
rect 24199 7590 24245 7642
rect 24269 7590 24315 7642
rect 24315 7590 24325 7642
rect 24349 7590 24379 7642
rect 24379 7590 24405 7642
rect 24109 7588 24165 7590
rect 24189 7588 24245 7590
rect 24269 7588 24325 7590
rect 24349 7588 24405 7590
rect 19478 7098 19534 7100
rect 19558 7098 19614 7100
rect 19638 7098 19694 7100
rect 19718 7098 19774 7100
rect 19478 7046 19504 7098
rect 19504 7046 19534 7098
rect 19558 7046 19568 7098
rect 19568 7046 19614 7098
rect 19638 7046 19684 7098
rect 19684 7046 19694 7098
rect 19718 7046 19748 7098
rect 19748 7046 19774 7098
rect 19478 7044 19534 7046
rect 19558 7044 19614 7046
rect 19638 7044 19694 7046
rect 19718 7044 19774 7046
rect 14848 6554 14904 6556
rect 14928 6554 14984 6556
rect 15008 6554 15064 6556
rect 15088 6554 15144 6556
rect 14848 6502 14874 6554
rect 14874 6502 14904 6554
rect 14928 6502 14938 6554
rect 14938 6502 14984 6554
rect 15008 6502 15054 6554
rect 15054 6502 15064 6554
rect 15088 6502 15118 6554
rect 15118 6502 15144 6554
rect 14848 6500 14904 6502
rect 14928 6500 14984 6502
rect 15008 6500 15064 6502
rect 15088 6500 15144 6502
rect 24109 6554 24165 6556
rect 24189 6554 24245 6556
rect 24269 6554 24325 6556
rect 24349 6554 24405 6556
rect 24109 6502 24135 6554
rect 24135 6502 24165 6554
rect 24189 6502 24199 6554
rect 24199 6502 24245 6554
rect 24269 6502 24315 6554
rect 24315 6502 24325 6554
rect 24349 6502 24379 6554
rect 24379 6502 24405 6554
rect 24109 6500 24165 6502
rect 24189 6500 24245 6502
rect 24269 6500 24325 6502
rect 24349 6500 24405 6502
rect 14848 5466 14904 5468
rect 14928 5466 14984 5468
rect 15008 5466 15064 5468
rect 15088 5466 15144 5468
rect 14848 5414 14874 5466
rect 14874 5414 14904 5466
rect 14928 5414 14938 5466
rect 14938 5414 14984 5466
rect 15008 5414 15054 5466
rect 15054 5414 15064 5466
rect 15088 5414 15118 5466
rect 15118 5414 15144 5466
rect 14848 5412 14904 5414
rect 14928 5412 14984 5414
rect 15008 5412 15064 5414
rect 15088 5412 15144 5414
rect 14848 4378 14904 4380
rect 14928 4378 14984 4380
rect 15008 4378 15064 4380
rect 15088 4378 15144 4380
rect 14848 4326 14874 4378
rect 14874 4326 14904 4378
rect 14928 4326 14938 4378
rect 14938 4326 14984 4378
rect 15008 4326 15054 4378
rect 15054 4326 15064 4378
rect 15088 4326 15118 4378
rect 15118 4326 15144 4378
rect 14848 4324 14904 4326
rect 14928 4324 14984 4326
rect 15008 4324 15064 4326
rect 15088 4324 15144 4326
rect 19478 6010 19534 6012
rect 19558 6010 19614 6012
rect 19638 6010 19694 6012
rect 19718 6010 19774 6012
rect 19478 5958 19504 6010
rect 19504 5958 19534 6010
rect 19558 5958 19568 6010
rect 19568 5958 19614 6010
rect 19638 5958 19684 6010
rect 19684 5958 19694 6010
rect 19718 5958 19748 6010
rect 19748 5958 19774 6010
rect 19478 5956 19534 5958
rect 19558 5956 19614 5958
rect 19638 5956 19694 5958
rect 19718 5956 19774 5958
rect 24109 5466 24165 5468
rect 24189 5466 24245 5468
rect 24269 5466 24325 5468
rect 24349 5466 24405 5468
rect 24109 5414 24135 5466
rect 24135 5414 24165 5466
rect 24189 5414 24199 5466
rect 24199 5414 24245 5466
rect 24269 5414 24315 5466
rect 24315 5414 24325 5466
rect 24349 5414 24379 5466
rect 24379 5414 24405 5466
rect 24109 5412 24165 5414
rect 24189 5412 24245 5414
rect 24269 5412 24325 5414
rect 24349 5412 24405 5414
rect 19478 4922 19534 4924
rect 19558 4922 19614 4924
rect 19638 4922 19694 4924
rect 19718 4922 19774 4924
rect 19478 4870 19504 4922
rect 19504 4870 19534 4922
rect 19558 4870 19568 4922
rect 19568 4870 19614 4922
rect 19638 4870 19684 4922
rect 19684 4870 19694 4922
rect 19718 4870 19748 4922
rect 19748 4870 19774 4922
rect 19478 4868 19534 4870
rect 19558 4868 19614 4870
rect 19638 4868 19694 4870
rect 19718 4868 19774 4870
rect 14848 3290 14904 3292
rect 14928 3290 14984 3292
rect 15008 3290 15064 3292
rect 15088 3290 15144 3292
rect 14848 3238 14874 3290
rect 14874 3238 14904 3290
rect 14928 3238 14938 3290
rect 14938 3238 14984 3290
rect 15008 3238 15054 3290
rect 15054 3238 15064 3290
rect 15088 3238 15118 3290
rect 15118 3238 15144 3290
rect 14848 3236 14904 3238
rect 14928 3236 14984 3238
rect 15008 3236 15064 3238
rect 15088 3236 15144 3238
rect 24109 4378 24165 4380
rect 24189 4378 24245 4380
rect 24269 4378 24325 4380
rect 24349 4378 24405 4380
rect 24109 4326 24135 4378
rect 24135 4326 24165 4378
rect 24189 4326 24199 4378
rect 24199 4326 24245 4378
rect 24269 4326 24315 4378
rect 24315 4326 24325 4378
rect 24349 4326 24379 4378
rect 24379 4326 24405 4378
rect 24109 4324 24165 4326
rect 24189 4324 24245 4326
rect 24269 4324 24325 4326
rect 24349 4324 24405 4326
rect 19478 3834 19534 3836
rect 19558 3834 19614 3836
rect 19638 3834 19694 3836
rect 19718 3834 19774 3836
rect 19478 3782 19504 3834
rect 19504 3782 19534 3834
rect 19558 3782 19568 3834
rect 19568 3782 19614 3834
rect 19638 3782 19684 3834
rect 19684 3782 19694 3834
rect 19718 3782 19748 3834
rect 19748 3782 19774 3834
rect 19478 3780 19534 3782
rect 19558 3780 19614 3782
rect 19638 3780 19694 3782
rect 19718 3780 19774 3782
rect 24109 3290 24165 3292
rect 24189 3290 24245 3292
rect 24269 3290 24325 3292
rect 24349 3290 24405 3292
rect 24109 3238 24135 3290
rect 24135 3238 24165 3290
rect 24189 3238 24199 3290
rect 24199 3238 24245 3290
rect 24269 3238 24315 3290
rect 24315 3238 24325 3290
rect 24349 3238 24379 3290
rect 24379 3238 24405 3290
rect 24109 3236 24165 3238
rect 24189 3236 24245 3238
rect 24269 3236 24325 3238
rect 24349 3236 24405 3238
rect 19478 2746 19534 2748
rect 19558 2746 19614 2748
rect 19638 2746 19694 2748
rect 19718 2746 19774 2748
rect 19478 2694 19504 2746
rect 19504 2694 19534 2746
rect 19558 2694 19568 2746
rect 19568 2694 19614 2746
rect 19638 2694 19684 2746
rect 19684 2694 19694 2746
rect 19718 2694 19748 2746
rect 19748 2694 19774 2746
rect 19478 2692 19534 2694
rect 19558 2692 19614 2694
rect 19638 2692 19694 2694
rect 19718 2692 19774 2694
rect 14848 2202 14904 2204
rect 14928 2202 14984 2204
rect 15008 2202 15064 2204
rect 15088 2202 15144 2204
rect 14848 2150 14874 2202
rect 14874 2150 14904 2202
rect 14928 2150 14938 2202
rect 14938 2150 14984 2202
rect 15008 2150 15054 2202
rect 15054 2150 15064 2202
rect 15088 2150 15118 2202
rect 15118 2150 15144 2202
rect 14848 2148 14904 2150
rect 14928 2148 14984 2150
rect 15008 2148 15064 2150
rect 15088 2148 15144 2150
rect 24109 2202 24165 2204
rect 24189 2202 24245 2204
rect 24269 2202 24325 2204
rect 24349 2202 24405 2204
rect 24109 2150 24135 2202
rect 24135 2150 24165 2202
rect 24189 2150 24199 2202
rect 24199 2150 24245 2202
rect 24269 2150 24315 2202
rect 24315 2150 24325 2202
rect 24349 2150 24379 2202
rect 24379 2150 24405 2202
rect 24109 2148 24165 2150
rect 24189 2148 24245 2150
rect 24269 2148 24325 2150
rect 24349 2148 24405 2150
rect 27158 2080 27214 2136
<< metal3 >>
rect 0 30018 800 30048
rect 1393 30018 1459 30021
rect 0 30016 1459 30018
rect 0 29960 1398 30016
rect 1454 29960 1459 30016
rect 0 29958 1459 29960
rect 0 29928 800 29958
rect 1393 29955 1459 29958
rect 10205 29952 10525 29953
rect 10205 29888 10213 29952
rect 10277 29888 10293 29952
rect 10357 29888 10373 29952
rect 10437 29888 10453 29952
rect 10517 29888 10525 29952
rect 10205 29887 10525 29888
rect 19466 29952 19786 29953
rect 19466 29888 19474 29952
rect 19538 29888 19554 29952
rect 19618 29888 19634 29952
rect 19698 29888 19714 29952
rect 19778 29888 19786 29952
rect 19466 29887 19786 29888
rect 5574 29408 5894 29409
rect 5574 29344 5582 29408
rect 5646 29344 5662 29408
rect 5726 29344 5742 29408
rect 5806 29344 5822 29408
rect 5886 29344 5894 29408
rect 5574 29343 5894 29344
rect 14836 29408 15156 29409
rect 14836 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15156 29408
rect 14836 29343 15156 29344
rect 24097 29408 24417 29409
rect 24097 29344 24105 29408
rect 24169 29344 24185 29408
rect 24249 29344 24265 29408
rect 24329 29344 24345 29408
rect 24409 29344 24417 29408
rect 24097 29343 24417 29344
rect 10205 28864 10525 28865
rect 10205 28800 10213 28864
rect 10277 28800 10293 28864
rect 10357 28800 10373 28864
rect 10437 28800 10453 28864
rect 10517 28800 10525 28864
rect 10205 28799 10525 28800
rect 19466 28864 19786 28865
rect 19466 28800 19474 28864
rect 19538 28800 19554 28864
rect 19618 28800 19634 28864
rect 19698 28800 19714 28864
rect 19778 28800 19786 28864
rect 19466 28799 19786 28800
rect 5574 28320 5894 28321
rect 5574 28256 5582 28320
rect 5646 28256 5662 28320
rect 5726 28256 5742 28320
rect 5806 28256 5822 28320
rect 5886 28256 5894 28320
rect 5574 28255 5894 28256
rect 14836 28320 15156 28321
rect 14836 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15156 28320
rect 14836 28255 15156 28256
rect 24097 28320 24417 28321
rect 24097 28256 24105 28320
rect 24169 28256 24185 28320
rect 24249 28256 24265 28320
rect 24329 28256 24345 28320
rect 24409 28256 24417 28320
rect 24097 28255 24417 28256
rect 10205 27776 10525 27777
rect 10205 27712 10213 27776
rect 10277 27712 10293 27776
rect 10357 27712 10373 27776
rect 10437 27712 10453 27776
rect 10517 27712 10525 27776
rect 10205 27711 10525 27712
rect 19466 27776 19786 27777
rect 19466 27712 19474 27776
rect 19538 27712 19554 27776
rect 19618 27712 19634 27776
rect 19698 27712 19714 27776
rect 19778 27712 19786 27776
rect 19466 27711 19786 27712
rect 5574 27232 5894 27233
rect 5574 27168 5582 27232
rect 5646 27168 5662 27232
rect 5726 27168 5742 27232
rect 5806 27168 5822 27232
rect 5886 27168 5894 27232
rect 5574 27167 5894 27168
rect 14836 27232 15156 27233
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 27167 15156 27168
rect 24097 27232 24417 27233
rect 24097 27168 24105 27232
rect 24169 27168 24185 27232
rect 24249 27168 24265 27232
rect 24329 27168 24345 27232
rect 24409 27168 24417 27232
rect 24097 27167 24417 27168
rect 10205 26688 10525 26689
rect 10205 26624 10213 26688
rect 10277 26624 10293 26688
rect 10357 26624 10373 26688
rect 10437 26624 10453 26688
rect 10517 26624 10525 26688
rect 10205 26623 10525 26624
rect 19466 26688 19786 26689
rect 19466 26624 19474 26688
rect 19538 26624 19554 26688
rect 19618 26624 19634 26688
rect 19698 26624 19714 26688
rect 19778 26624 19786 26688
rect 19466 26623 19786 26624
rect 5574 26144 5894 26145
rect 5574 26080 5582 26144
rect 5646 26080 5662 26144
rect 5726 26080 5742 26144
rect 5806 26080 5822 26144
rect 5886 26080 5894 26144
rect 5574 26079 5894 26080
rect 14836 26144 15156 26145
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 26079 15156 26080
rect 24097 26144 24417 26145
rect 24097 26080 24105 26144
rect 24169 26080 24185 26144
rect 24249 26080 24265 26144
rect 24329 26080 24345 26144
rect 24409 26080 24417 26144
rect 24097 26079 24417 26080
rect 10205 25600 10525 25601
rect 10205 25536 10213 25600
rect 10277 25536 10293 25600
rect 10357 25536 10373 25600
rect 10437 25536 10453 25600
rect 10517 25536 10525 25600
rect 10205 25535 10525 25536
rect 19466 25600 19786 25601
rect 19466 25536 19474 25600
rect 19538 25536 19554 25600
rect 19618 25536 19634 25600
rect 19698 25536 19714 25600
rect 19778 25536 19786 25600
rect 19466 25535 19786 25536
rect 5574 25056 5894 25057
rect 5574 24992 5582 25056
rect 5646 24992 5662 25056
rect 5726 24992 5742 25056
rect 5806 24992 5822 25056
rect 5886 24992 5894 25056
rect 5574 24991 5894 24992
rect 14836 25056 15156 25057
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 24991 15156 24992
rect 24097 25056 24417 25057
rect 24097 24992 24105 25056
rect 24169 24992 24185 25056
rect 24249 24992 24265 25056
rect 24329 24992 24345 25056
rect 24409 24992 24417 25056
rect 24097 24991 24417 24992
rect 10205 24512 10525 24513
rect 10205 24448 10213 24512
rect 10277 24448 10293 24512
rect 10357 24448 10373 24512
rect 10437 24448 10453 24512
rect 10517 24448 10525 24512
rect 10205 24447 10525 24448
rect 19466 24512 19786 24513
rect 19466 24448 19474 24512
rect 19538 24448 19554 24512
rect 19618 24448 19634 24512
rect 19698 24448 19714 24512
rect 19778 24448 19786 24512
rect 19466 24447 19786 24448
rect 5574 23968 5894 23969
rect 5574 23904 5582 23968
rect 5646 23904 5662 23968
rect 5726 23904 5742 23968
rect 5806 23904 5822 23968
rect 5886 23904 5894 23968
rect 5574 23903 5894 23904
rect 14836 23968 15156 23969
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 23903 15156 23904
rect 24097 23968 24417 23969
rect 24097 23904 24105 23968
rect 24169 23904 24185 23968
rect 24249 23904 24265 23968
rect 24329 23904 24345 23968
rect 24409 23904 24417 23968
rect 24097 23903 24417 23904
rect 10205 23424 10525 23425
rect 10205 23360 10213 23424
rect 10277 23360 10293 23424
rect 10357 23360 10373 23424
rect 10437 23360 10453 23424
rect 10517 23360 10525 23424
rect 10205 23359 10525 23360
rect 19466 23424 19786 23425
rect 19466 23360 19474 23424
rect 19538 23360 19554 23424
rect 19618 23360 19634 23424
rect 19698 23360 19714 23424
rect 19778 23360 19786 23424
rect 19466 23359 19786 23360
rect 5574 22880 5894 22881
rect 5574 22816 5582 22880
rect 5646 22816 5662 22880
rect 5726 22816 5742 22880
rect 5806 22816 5822 22880
rect 5886 22816 5894 22880
rect 5574 22815 5894 22816
rect 14836 22880 15156 22881
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 22815 15156 22816
rect 24097 22880 24417 22881
rect 24097 22816 24105 22880
rect 24169 22816 24185 22880
rect 24249 22816 24265 22880
rect 24329 22816 24345 22880
rect 24409 22816 24417 22880
rect 24097 22815 24417 22816
rect 10205 22336 10525 22337
rect 10205 22272 10213 22336
rect 10277 22272 10293 22336
rect 10357 22272 10373 22336
rect 10437 22272 10453 22336
rect 10517 22272 10525 22336
rect 10205 22271 10525 22272
rect 19466 22336 19786 22337
rect 19466 22272 19474 22336
rect 19538 22272 19554 22336
rect 19618 22272 19634 22336
rect 19698 22272 19714 22336
rect 19778 22272 19786 22336
rect 19466 22271 19786 22272
rect 5574 21792 5894 21793
rect 5574 21728 5582 21792
rect 5646 21728 5662 21792
rect 5726 21728 5742 21792
rect 5806 21728 5822 21792
rect 5886 21728 5894 21792
rect 5574 21727 5894 21728
rect 14836 21792 15156 21793
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 21727 15156 21728
rect 24097 21792 24417 21793
rect 24097 21728 24105 21792
rect 24169 21728 24185 21792
rect 24249 21728 24265 21792
rect 24329 21728 24345 21792
rect 24409 21728 24417 21792
rect 24097 21727 24417 21728
rect 10205 21248 10525 21249
rect 10205 21184 10213 21248
rect 10277 21184 10293 21248
rect 10357 21184 10373 21248
rect 10437 21184 10453 21248
rect 10517 21184 10525 21248
rect 10205 21183 10525 21184
rect 19466 21248 19786 21249
rect 19466 21184 19474 21248
rect 19538 21184 19554 21248
rect 19618 21184 19634 21248
rect 19698 21184 19714 21248
rect 19778 21184 19786 21248
rect 19466 21183 19786 21184
rect 5574 20704 5894 20705
rect 5574 20640 5582 20704
rect 5646 20640 5662 20704
rect 5726 20640 5742 20704
rect 5806 20640 5822 20704
rect 5886 20640 5894 20704
rect 5574 20639 5894 20640
rect 14836 20704 15156 20705
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 20639 15156 20640
rect 24097 20704 24417 20705
rect 24097 20640 24105 20704
rect 24169 20640 24185 20704
rect 24249 20640 24265 20704
rect 24329 20640 24345 20704
rect 24409 20640 24417 20704
rect 24097 20639 24417 20640
rect 10205 20160 10525 20161
rect 10205 20096 10213 20160
rect 10277 20096 10293 20160
rect 10357 20096 10373 20160
rect 10437 20096 10453 20160
rect 10517 20096 10525 20160
rect 10205 20095 10525 20096
rect 19466 20160 19786 20161
rect 19466 20096 19474 20160
rect 19538 20096 19554 20160
rect 19618 20096 19634 20160
rect 19698 20096 19714 20160
rect 19778 20096 19786 20160
rect 19466 20095 19786 20096
rect 5574 19616 5894 19617
rect 5574 19552 5582 19616
rect 5646 19552 5662 19616
rect 5726 19552 5742 19616
rect 5806 19552 5822 19616
rect 5886 19552 5894 19616
rect 5574 19551 5894 19552
rect 14836 19616 15156 19617
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 19551 15156 19552
rect 24097 19616 24417 19617
rect 24097 19552 24105 19616
rect 24169 19552 24185 19616
rect 24249 19552 24265 19616
rect 24329 19552 24345 19616
rect 24409 19552 24417 19616
rect 24097 19551 24417 19552
rect 10205 19072 10525 19073
rect 10205 19008 10213 19072
rect 10277 19008 10293 19072
rect 10357 19008 10373 19072
rect 10437 19008 10453 19072
rect 10517 19008 10525 19072
rect 10205 19007 10525 19008
rect 19466 19072 19786 19073
rect 19466 19008 19474 19072
rect 19538 19008 19554 19072
rect 19618 19008 19634 19072
rect 19698 19008 19714 19072
rect 19778 19008 19786 19072
rect 19466 19007 19786 19008
rect 5574 18528 5894 18529
rect 5574 18464 5582 18528
rect 5646 18464 5662 18528
rect 5726 18464 5742 18528
rect 5806 18464 5822 18528
rect 5886 18464 5894 18528
rect 5574 18463 5894 18464
rect 14836 18528 15156 18529
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 18463 15156 18464
rect 24097 18528 24417 18529
rect 24097 18464 24105 18528
rect 24169 18464 24185 18528
rect 24249 18464 24265 18528
rect 24329 18464 24345 18528
rect 24409 18464 24417 18528
rect 24097 18463 24417 18464
rect 10205 17984 10525 17985
rect 10205 17920 10213 17984
rect 10277 17920 10293 17984
rect 10357 17920 10373 17984
rect 10437 17920 10453 17984
rect 10517 17920 10525 17984
rect 10205 17919 10525 17920
rect 19466 17984 19786 17985
rect 19466 17920 19474 17984
rect 19538 17920 19554 17984
rect 19618 17920 19634 17984
rect 19698 17920 19714 17984
rect 19778 17920 19786 17984
rect 19466 17919 19786 17920
rect 5574 17440 5894 17441
rect 5574 17376 5582 17440
rect 5646 17376 5662 17440
rect 5726 17376 5742 17440
rect 5806 17376 5822 17440
rect 5886 17376 5894 17440
rect 5574 17375 5894 17376
rect 14836 17440 15156 17441
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 17375 15156 17376
rect 24097 17440 24417 17441
rect 24097 17376 24105 17440
rect 24169 17376 24185 17440
rect 24249 17376 24265 17440
rect 24329 17376 24345 17440
rect 24409 17376 24417 17440
rect 24097 17375 24417 17376
rect 28165 17098 28231 17101
rect 29224 17098 30024 17128
rect 28165 17096 30024 17098
rect 28165 17040 28170 17096
rect 28226 17040 30024 17096
rect 28165 17038 30024 17040
rect 28165 17035 28231 17038
rect 29224 17008 30024 17038
rect 10205 16896 10525 16897
rect 10205 16832 10213 16896
rect 10277 16832 10293 16896
rect 10357 16832 10373 16896
rect 10437 16832 10453 16896
rect 10517 16832 10525 16896
rect 10205 16831 10525 16832
rect 19466 16896 19786 16897
rect 19466 16832 19474 16896
rect 19538 16832 19554 16896
rect 19618 16832 19634 16896
rect 19698 16832 19714 16896
rect 19778 16832 19786 16896
rect 19466 16831 19786 16832
rect 5574 16352 5894 16353
rect 5574 16288 5582 16352
rect 5646 16288 5662 16352
rect 5726 16288 5742 16352
rect 5806 16288 5822 16352
rect 5886 16288 5894 16352
rect 5574 16287 5894 16288
rect 14836 16352 15156 16353
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 16287 15156 16288
rect 24097 16352 24417 16353
rect 24097 16288 24105 16352
rect 24169 16288 24185 16352
rect 24249 16288 24265 16352
rect 24329 16288 24345 16352
rect 24409 16288 24417 16352
rect 24097 16287 24417 16288
rect 10205 15808 10525 15809
rect 10205 15744 10213 15808
rect 10277 15744 10293 15808
rect 10357 15744 10373 15808
rect 10437 15744 10453 15808
rect 10517 15744 10525 15808
rect 10205 15743 10525 15744
rect 19466 15808 19786 15809
rect 19466 15744 19474 15808
rect 19538 15744 19554 15808
rect 19618 15744 19634 15808
rect 19698 15744 19714 15808
rect 19778 15744 19786 15808
rect 19466 15743 19786 15744
rect 5574 15264 5894 15265
rect 5574 15200 5582 15264
rect 5646 15200 5662 15264
rect 5726 15200 5742 15264
rect 5806 15200 5822 15264
rect 5886 15200 5894 15264
rect 5574 15199 5894 15200
rect 14836 15264 15156 15265
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 15199 15156 15200
rect 24097 15264 24417 15265
rect 24097 15200 24105 15264
rect 24169 15200 24185 15264
rect 24249 15200 24265 15264
rect 24329 15200 24345 15264
rect 24409 15200 24417 15264
rect 24097 15199 24417 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 10205 14720 10525 14721
rect 10205 14656 10213 14720
rect 10277 14656 10293 14720
rect 10357 14656 10373 14720
rect 10437 14656 10453 14720
rect 10517 14656 10525 14720
rect 10205 14655 10525 14656
rect 19466 14720 19786 14721
rect 19466 14656 19474 14720
rect 19538 14656 19554 14720
rect 19618 14656 19634 14720
rect 19698 14656 19714 14720
rect 19778 14656 19786 14720
rect 19466 14655 19786 14656
rect 5574 14176 5894 14177
rect 5574 14112 5582 14176
rect 5646 14112 5662 14176
rect 5726 14112 5742 14176
rect 5806 14112 5822 14176
rect 5886 14112 5894 14176
rect 5574 14111 5894 14112
rect 14836 14176 15156 14177
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 14111 15156 14112
rect 24097 14176 24417 14177
rect 24097 14112 24105 14176
rect 24169 14112 24185 14176
rect 24249 14112 24265 14176
rect 24329 14112 24345 14176
rect 24409 14112 24417 14176
rect 24097 14111 24417 14112
rect 10205 13632 10525 13633
rect 10205 13568 10213 13632
rect 10277 13568 10293 13632
rect 10357 13568 10373 13632
rect 10437 13568 10453 13632
rect 10517 13568 10525 13632
rect 10205 13567 10525 13568
rect 19466 13632 19786 13633
rect 19466 13568 19474 13632
rect 19538 13568 19554 13632
rect 19618 13568 19634 13632
rect 19698 13568 19714 13632
rect 19778 13568 19786 13632
rect 19466 13567 19786 13568
rect 5574 13088 5894 13089
rect 5574 13024 5582 13088
rect 5646 13024 5662 13088
rect 5726 13024 5742 13088
rect 5806 13024 5822 13088
rect 5886 13024 5894 13088
rect 5574 13023 5894 13024
rect 14836 13088 15156 13089
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 13023 15156 13024
rect 24097 13088 24417 13089
rect 24097 13024 24105 13088
rect 24169 13024 24185 13088
rect 24249 13024 24265 13088
rect 24329 13024 24345 13088
rect 24409 13024 24417 13088
rect 24097 13023 24417 13024
rect 10205 12544 10525 12545
rect 10205 12480 10213 12544
rect 10277 12480 10293 12544
rect 10357 12480 10373 12544
rect 10437 12480 10453 12544
rect 10517 12480 10525 12544
rect 10205 12479 10525 12480
rect 19466 12544 19786 12545
rect 19466 12480 19474 12544
rect 19538 12480 19554 12544
rect 19618 12480 19634 12544
rect 19698 12480 19714 12544
rect 19778 12480 19786 12544
rect 19466 12479 19786 12480
rect 5574 12000 5894 12001
rect 5574 11936 5582 12000
rect 5646 11936 5662 12000
rect 5726 11936 5742 12000
rect 5806 11936 5822 12000
rect 5886 11936 5894 12000
rect 5574 11935 5894 11936
rect 14836 12000 15156 12001
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 11935 15156 11936
rect 24097 12000 24417 12001
rect 24097 11936 24105 12000
rect 24169 11936 24185 12000
rect 24249 11936 24265 12000
rect 24329 11936 24345 12000
rect 24409 11936 24417 12000
rect 24097 11935 24417 11936
rect 10205 11456 10525 11457
rect 10205 11392 10213 11456
rect 10277 11392 10293 11456
rect 10357 11392 10373 11456
rect 10437 11392 10453 11456
rect 10517 11392 10525 11456
rect 10205 11391 10525 11392
rect 19466 11456 19786 11457
rect 19466 11392 19474 11456
rect 19538 11392 19554 11456
rect 19618 11392 19634 11456
rect 19698 11392 19714 11456
rect 19778 11392 19786 11456
rect 19466 11391 19786 11392
rect 5574 10912 5894 10913
rect 5574 10848 5582 10912
rect 5646 10848 5662 10912
rect 5726 10848 5742 10912
rect 5806 10848 5822 10912
rect 5886 10848 5894 10912
rect 5574 10847 5894 10848
rect 14836 10912 15156 10913
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 10847 15156 10848
rect 24097 10912 24417 10913
rect 24097 10848 24105 10912
rect 24169 10848 24185 10912
rect 24249 10848 24265 10912
rect 24329 10848 24345 10912
rect 24409 10848 24417 10912
rect 24097 10847 24417 10848
rect 10205 10368 10525 10369
rect 10205 10304 10213 10368
rect 10277 10304 10293 10368
rect 10357 10304 10373 10368
rect 10437 10304 10453 10368
rect 10517 10304 10525 10368
rect 10205 10303 10525 10304
rect 19466 10368 19786 10369
rect 19466 10304 19474 10368
rect 19538 10304 19554 10368
rect 19618 10304 19634 10368
rect 19698 10304 19714 10368
rect 19778 10304 19786 10368
rect 19466 10303 19786 10304
rect 5574 9824 5894 9825
rect 5574 9760 5582 9824
rect 5646 9760 5662 9824
rect 5726 9760 5742 9824
rect 5806 9760 5822 9824
rect 5886 9760 5894 9824
rect 5574 9759 5894 9760
rect 14836 9824 15156 9825
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 9759 15156 9760
rect 24097 9824 24417 9825
rect 24097 9760 24105 9824
rect 24169 9760 24185 9824
rect 24249 9760 24265 9824
rect 24329 9760 24345 9824
rect 24409 9760 24417 9824
rect 24097 9759 24417 9760
rect 10205 9280 10525 9281
rect 10205 9216 10213 9280
rect 10277 9216 10293 9280
rect 10357 9216 10373 9280
rect 10437 9216 10453 9280
rect 10517 9216 10525 9280
rect 10205 9215 10525 9216
rect 19466 9280 19786 9281
rect 19466 9216 19474 9280
rect 19538 9216 19554 9280
rect 19618 9216 19634 9280
rect 19698 9216 19714 9280
rect 19778 9216 19786 9280
rect 19466 9215 19786 9216
rect 5574 8736 5894 8737
rect 5574 8672 5582 8736
rect 5646 8672 5662 8736
rect 5726 8672 5742 8736
rect 5806 8672 5822 8736
rect 5886 8672 5894 8736
rect 5574 8671 5894 8672
rect 14836 8736 15156 8737
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 8671 15156 8672
rect 24097 8736 24417 8737
rect 24097 8672 24105 8736
rect 24169 8672 24185 8736
rect 24249 8672 24265 8736
rect 24329 8672 24345 8736
rect 24409 8672 24417 8736
rect 24097 8671 24417 8672
rect 10205 8192 10525 8193
rect 10205 8128 10213 8192
rect 10277 8128 10293 8192
rect 10357 8128 10373 8192
rect 10437 8128 10453 8192
rect 10517 8128 10525 8192
rect 10205 8127 10525 8128
rect 19466 8192 19786 8193
rect 19466 8128 19474 8192
rect 19538 8128 19554 8192
rect 19618 8128 19634 8192
rect 19698 8128 19714 8192
rect 19778 8128 19786 8192
rect 19466 8127 19786 8128
rect 5574 7648 5894 7649
rect 5574 7584 5582 7648
rect 5646 7584 5662 7648
rect 5726 7584 5742 7648
rect 5806 7584 5822 7648
rect 5886 7584 5894 7648
rect 5574 7583 5894 7584
rect 14836 7648 15156 7649
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 7583 15156 7584
rect 24097 7648 24417 7649
rect 24097 7584 24105 7648
rect 24169 7584 24185 7648
rect 24249 7584 24265 7648
rect 24329 7584 24345 7648
rect 24409 7584 24417 7648
rect 24097 7583 24417 7584
rect 10205 7104 10525 7105
rect 10205 7040 10213 7104
rect 10277 7040 10293 7104
rect 10357 7040 10373 7104
rect 10437 7040 10453 7104
rect 10517 7040 10525 7104
rect 10205 7039 10525 7040
rect 19466 7104 19786 7105
rect 19466 7040 19474 7104
rect 19538 7040 19554 7104
rect 19618 7040 19634 7104
rect 19698 7040 19714 7104
rect 19778 7040 19786 7104
rect 19466 7039 19786 7040
rect 5574 6560 5894 6561
rect 5574 6496 5582 6560
rect 5646 6496 5662 6560
rect 5726 6496 5742 6560
rect 5806 6496 5822 6560
rect 5886 6496 5894 6560
rect 5574 6495 5894 6496
rect 14836 6560 15156 6561
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 6495 15156 6496
rect 24097 6560 24417 6561
rect 24097 6496 24105 6560
rect 24169 6496 24185 6560
rect 24249 6496 24265 6560
rect 24329 6496 24345 6560
rect 24409 6496 24417 6560
rect 24097 6495 24417 6496
rect 10205 6016 10525 6017
rect 10205 5952 10213 6016
rect 10277 5952 10293 6016
rect 10357 5952 10373 6016
rect 10437 5952 10453 6016
rect 10517 5952 10525 6016
rect 10205 5951 10525 5952
rect 19466 6016 19786 6017
rect 19466 5952 19474 6016
rect 19538 5952 19554 6016
rect 19618 5952 19634 6016
rect 19698 5952 19714 6016
rect 19778 5952 19786 6016
rect 19466 5951 19786 5952
rect 5574 5472 5894 5473
rect 5574 5408 5582 5472
rect 5646 5408 5662 5472
rect 5726 5408 5742 5472
rect 5806 5408 5822 5472
rect 5886 5408 5894 5472
rect 5574 5407 5894 5408
rect 14836 5472 15156 5473
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 5407 15156 5408
rect 24097 5472 24417 5473
rect 24097 5408 24105 5472
rect 24169 5408 24185 5472
rect 24249 5408 24265 5472
rect 24329 5408 24345 5472
rect 24409 5408 24417 5472
rect 24097 5407 24417 5408
rect 10205 4928 10525 4929
rect 10205 4864 10213 4928
rect 10277 4864 10293 4928
rect 10357 4864 10373 4928
rect 10437 4864 10453 4928
rect 10517 4864 10525 4928
rect 10205 4863 10525 4864
rect 19466 4928 19786 4929
rect 19466 4864 19474 4928
rect 19538 4864 19554 4928
rect 19618 4864 19634 4928
rect 19698 4864 19714 4928
rect 19778 4864 19786 4928
rect 19466 4863 19786 4864
rect 5574 4384 5894 4385
rect 5574 4320 5582 4384
rect 5646 4320 5662 4384
rect 5726 4320 5742 4384
rect 5806 4320 5822 4384
rect 5886 4320 5894 4384
rect 5574 4319 5894 4320
rect 14836 4384 15156 4385
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 4319 15156 4320
rect 24097 4384 24417 4385
rect 24097 4320 24105 4384
rect 24169 4320 24185 4384
rect 24249 4320 24265 4384
rect 24329 4320 24345 4384
rect 24409 4320 24417 4384
rect 24097 4319 24417 4320
rect 10205 3840 10525 3841
rect 10205 3776 10213 3840
rect 10277 3776 10293 3840
rect 10357 3776 10373 3840
rect 10437 3776 10453 3840
rect 10517 3776 10525 3840
rect 10205 3775 10525 3776
rect 19466 3840 19786 3841
rect 19466 3776 19474 3840
rect 19538 3776 19554 3840
rect 19618 3776 19634 3840
rect 19698 3776 19714 3840
rect 19778 3776 19786 3840
rect 19466 3775 19786 3776
rect 5574 3296 5894 3297
rect 5574 3232 5582 3296
rect 5646 3232 5662 3296
rect 5726 3232 5742 3296
rect 5806 3232 5822 3296
rect 5886 3232 5894 3296
rect 5574 3231 5894 3232
rect 14836 3296 15156 3297
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 3231 15156 3232
rect 24097 3296 24417 3297
rect 24097 3232 24105 3296
rect 24169 3232 24185 3296
rect 24249 3232 24265 3296
rect 24329 3232 24345 3296
rect 24409 3232 24417 3296
rect 24097 3231 24417 3232
rect 10205 2752 10525 2753
rect 10205 2688 10213 2752
rect 10277 2688 10293 2752
rect 10357 2688 10373 2752
rect 10437 2688 10453 2752
rect 10517 2688 10525 2752
rect 10205 2687 10525 2688
rect 19466 2752 19786 2753
rect 19466 2688 19474 2752
rect 19538 2688 19554 2752
rect 19618 2688 19634 2752
rect 19698 2688 19714 2752
rect 19778 2688 19786 2752
rect 19466 2687 19786 2688
rect 5574 2208 5894 2209
rect 5574 2144 5582 2208
rect 5646 2144 5662 2208
rect 5726 2144 5742 2208
rect 5806 2144 5822 2208
rect 5886 2144 5894 2208
rect 5574 2143 5894 2144
rect 14836 2208 15156 2209
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2143 15156 2144
rect 24097 2208 24417 2209
rect 24097 2144 24105 2208
rect 24169 2144 24185 2208
rect 24249 2144 24265 2208
rect 24329 2144 24345 2208
rect 24409 2144 24417 2208
rect 24097 2143 24417 2144
rect 27153 2138 27219 2141
rect 29224 2138 30024 2168
rect 27153 2136 30024 2138
rect 27153 2080 27158 2136
rect 27214 2080 30024 2136
rect 27153 2078 30024 2080
rect 27153 2075 27219 2078
rect 29224 2048 30024 2078
<< via3 >>
rect 10213 29948 10277 29952
rect 10213 29892 10217 29948
rect 10217 29892 10273 29948
rect 10273 29892 10277 29948
rect 10213 29888 10277 29892
rect 10293 29948 10357 29952
rect 10293 29892 10297 29948
rect 10297 29892 10353 29948
rect 10353 29892 10357 29948
rect 10293 29888 10357 29892
rect 10373 29948 10437 29952
rect 10373 29892 10377 29948
rect 10377 29892 10433 29948
rect 10433 29892 10437 29948
rect 10373 29888 10437 29892
rect 10453 29948 10517 29952
rect 10453 29892 10457 29948
rect 10457 29892 10513 29948
rect 10513 29892 10517 29948
rect 10453 29888 10517 29892
rect 19474 29948 19538 29952
rect 19474 29892 19478 29948
rect 19478 29892 19534 29948
rect 19534 29892 19538 29948
rect 19474 29888 19538 29892
rect 19554 29948 19618 29952
rect 19554 29892 19558 29948
rect 19558 29892 19614 29948
rect 19614 29892 19618 29948
rect 19554 29888 19618 29892
rect 19634 29948 19698 29952
rect 19634 29892 19638 29948
rect 19638 29892 19694 29948
rect 19694 29892 19698 29948
rect 19634 29888 19698 29892
rect 19714 29948 19778 29952
rect 19714 29892 19718 29948
rect 19718 29892 19774 29948
rect 19774 29892 19778 29948
rect 19714 29888 19778 29892
rect 5582 29404 5646 29408
rect 5582 29348 5586 29404
rect 5586 29348 5642 29404
rect 5642 29348 5646 29404
rect 5582 29344 5646 29348
rect 5662 29404 5726 29408
rect 5662 29348 5666 29404
rect 5666 29348 5722 29404
rect 5722 29348 5726 29404
rect 5662 29344 5726 29348
rect 5742 29404 5806 29408
rect 5742 29348 5746 29404
rect 5746 29348 5802 29404
rect 5802 29348 5806 29404
rect 5742 29344 5806 29348
rect 5822 29404 5886 29408
rect 5822 29348 5826 29404
rect 5826 29348 5882 29404
rect 5882 29348 5886 29404
rect 5822 29344 5886 29348
rect 14844 29404 14908 29408
rect 14844 29348 14848 29404
rect 14848 29348 14904 29404
rect 14904 29348 14908 29404
rect 14844 29344 14908 29348
rect 14924 29404 14988 29408
rect 14924 29348 14928 29404
rect 14928 29348 14984 29404
rect 14984 29348 14988 29404
rect 14924 29344 14988 29348
rect 15004 29404 15068 29408
rect 15004 29348 15008 29404
rect 15008 29348 15064 29404
rect 15064 29348 15068 29404
rect 15004 29344 15068 29348
rect 15084 29404 15148 29408
rect 15084 29348 15088 29404
rect 15088 29348 15144 29404
rect 15144 29348 15148 29404
rect 15084 29344 15148 29348
rect 24105 29404 24169 29408
rect 24105 29348 24109 29404
rect 24109 29348 24165 29404
rect 24165 29348 24169 29404
rect 24105 29344 24169 29348
rect 24185 29404 24249 29408
rect 24185 29348 24189 29404
rect 24189 29348 24245 29404
rect 24245 29348 24249 29404
rect 24185 29344 24249 29348
rect 24265 29404 24329 29408
rect 24265 29348 24269 29404
rect 24269 29348 24325 29404
rect 24325 29348 24329 29404
rect 24265 29344 24329 29348
rect 24345 29404 24409 29408
rect 24345 29348 24349 29404
rect 24349 29348 24405 29404
rect 24405 29348 24409 29404
rect 24345 29344 24409 29348
rect 10213 28860 10277 28864
rect 10213 28804 10217 28860
rect 10217 28804 10273 28860
rect 10273 28804 10277 28860
rect 10213 28800 10277 28804
rect 10293 28860 10357 28864
rect 10293 28804 10297 28860
rect 10297 28804 10353 28860
rect 10353 28804 10357 28860
rect 10293 28800 10357 28804
rect 10373 28860 10437 28864
rect 10373 28804 10377 28860
rect 10377 28804 10433 28860
rect 10433 28804 10437 28860
rect 10373 28800 10437 28804
rect 10453 28860 10517 28864
rect 10453 28804 10457 28860
rect 10457 28804 10513 28860
rect 10513 28804 10517 28860
rect 10453 28800 10517 28804
rect 19474 28860 19538 28864
rect 19474 28804 19478 28860
rect 19478 28804 19534 28860
rect 19534 28804 19538 28860
rect 19474 28800 19538 28804
rect 19554 28860 19618 28864
rect 19554 28804 19558 28860
rect 19558 28804 19614 28860
rect 19614 28804 19618 28860
rect 19554 28800 19618 28804
rect 19634 28860 19698 28864
rect 19634 28804 19638 28860
rect 19638 28804 19694 28860
rect 19694 28804 19698 28860
rect 19634 28800 19698 28804
rect 19714 28860 19778 28864
rect 19714 28804 19718 28860
rect 19718 28804 19774 28860
rect 19774 28804 19778 28860
rect 19714 28800 19778 28804
rect 5582 28316 5646 28320
rect 5582 28260 5586 28316
rect 5586 28260 5642 28316
rect 5642 28260 5646 28316
rect 5582 28256 5646 28260
rect 5662 28316 5726 28320
rect 5662 28260 5666 28316
rect 5666 28260 5722 28316
rect 5722 28260 5726 28316
rect 5662 28256 5726 28260
rect 5742 28316 5806 28320
rect 5742 28260 5746 28316
rect 5746 28260 5802 28316
rect 5802 28260 5806 28316
rect 5742 28256 5806 28260
rect 5822 28316 5886 28320
rect 5822 28260 5826 28316
rect 5826 28260 5882 28316
rect 5882 28260 5886 28316
rect 5822 28256 5886 28260
rect 14844 28316 14908 28320
rect 14844 28260 14848 28316
rect 14848 28260 14904 28316
rect 14904 28260 14908 28316
rect 14844 28256 14908 28260
rect 14924 28316 14988 28320
rect 14924 28260 14928 28316
rect 14928 28260 14984 28316
rect 14984 28260 14988 28316
rect 14924 28256 14988 28260
rect 15004 28316 15068 28320
rect 15004 28260 15008 28316
rect 15008 28260 15064 28316
rect 15064 28260 15068 28316
rect 15004 28256 15068 28260
rect 15084 28316 15148 28320
rect 15084 28260 15088 28316
rect 15088 28260 15144 28316
rect 15144 28260 15148 28316
rect 15084 28256 15148 28260
rect 24105 28316 24169 28320
rect 24105 28260 24109 28316
rect 24109 28260 24165 28316
rect 24165 28260 24169 28316
rect 24105 28256 24169 28260
rect 24185 28316 24249 28320
rect 24185 28260 24189 28316
rect 24189 28260 24245 28316
rect 24245 28260 24249 28316
rect 24185 28256 24249 28260
rect 24265 28316 24329 28320
rect 24265 28260 24269 28316
rect 24269 28260 24325 28316
rect 24325 28260 24329 28316
rect 24265 28256 24329 28260
rect 24345 28316 24409 28320
rect 24345 28260 24349 28316
rect 24349 28260 24405 28316
rect 24405 28260 24409 28316
rect 24345 28256 24409 28260
rect 10213 27772 10277 27776
rect 10213 27716 10217 27772
rect 10217 27716 10273 27772
rect 10273 27716 10277 27772
rect 10213 27712 10277 27716
rect 10293 27772 10357 27776
rect 10293 27716 10297 27772
rect 10297 27716 10353 27772
rect 10353 27716 10357 27772
rect 10293 27712 10357 27716
rect 10373 27772 10437 27776
rect 10373 27716 10377 27772
rect 10377 27716 10433 27772
rect 10433 27716 10437 27772
rect 10373 27712 10437 27716
rect 10453 27772 10517 27776
rect 10453 27716 10457 27772
rect 10457 27716 10513 27772
rect 10513 27716 10517 27772
rect 10453 27712 10517 27716
rect 19474 27772 19538 27776
rect 19474 27716 19478 27772
rect 19478 27716 19534 27772
rect 19534 27716 19538 27772
rect 19474 27712 19538 27716
rect 19554 27772 19618 27776
rect 19554 27716 19558 27772
rect 19558 27716 19614 27772
rect 19614 27716 19618 27772
rect 19554 27712 19618 27716
rect 19634 27772 19698 27776
rect 19634 27716 19638 27772
rect 19638 27716 19694 27772
rect 19694 27716 19698 27772
rect 19634 27712 19698 27716
rect 19714 27772 19778 27776
rect 19714 27716 19718 27772
rect 19718 27716 19774 27772
rect 19774 27716 19778 27772
rect 19714 27712 19778 27716
rect 5582 27228 5646 27232
rect 5582 27172 5586 27228
rect 5586 27172 5642 27228
rect 5642 27172 5646 27228
rect 5582 27168 5646 27172
rect 5662 27228 5726 27232
rect 5662 27172 5666 27228
rect 5666 27172 5722 27228
rect 5722 27172 5726 27228
rect 5662 27168 5726 27172
rect 5742 27228 5806 27232
rect 5742 27172 5746 27228
rect 5746 27172 5802 27228
rect 5802 27172 5806 27228
rect 5742 27168 5806 27172
rect 5822 27228 5886 27232
rect 5822 27172 5826 27228
rect 5826 27172 5882 27228
rect 5882 27172 5886 27228
rect 5822 27168 5886 27172
rect 14844 27228 14908 27232
rect 14844 27172 14848 27228
rect 14848 27172 14904 27228
rect 14904 27172 14908 27228
rect 14844 27168 14908 27172
rect 14924 27228 14988 27232
rect 14924 27172 14928 27228
rect 14928 27172 14984 27228
rect 14984 27172 14988 27228
rect 14924 27168 14988 27172
rect 15004 27228 15068 27232
rect 15004 27172 15008 27228
rect 15008 27172 15064 27228
rect 15064 27172 15068 27228
rect 15004 27168 15068 27172
rect 15084 27228 15148 27232
rect 15084 27172 15088 27228
rect 15088 27172 15144 27228
rect 15144 27172 15148 27228
rect 15084 27168 15148 27172
rect 24105 27228 24169 27232
rect 24105 27172 24109 27228
rect 24109 27172 24165 27228
rect 24165 27172 24169 27228
rect 24105 27168 24169 27172
rect 24185 27228 24249 27232
rect 24185 27172 24189 27228
rect 24189 27172 24245 27228
rect 24245 27172 24249 27228
rect 24185 27168 24249 27172
rect 24265 27228 24329 27232
rect 24265 27172 24269 27228
rect 24269 27172 24325 27228
rect 24325 27172 24329 27228
rect 24265 27168 24329 27172
rect 24345 27228 24409 27232
rect 24345 27172 24349 27228
rect 24349 27172 24405 27228
rect 24405 27172 24409 27228
rect 24345 27168 24409 27172
rect 10213 26684 10277 26688
rect 10213 26628 10217 26684
rect 10217 26628 10273 26684
rect 10273 26628 10277 26684
rect 10213 26624 10277 26628
rect 10293 26684 10357 26688
rect 10293 26628 10297 26684
rect 10297 26628 10353 26684
rect 10353 26628 10357 26684
rect 10293 26624 10357 26628
rect 10373 26684 10437 26688
rect 10373 26628 10377 26684
rect 10377 26628 10433 26684
rect 10433 26628 10437 26684
rect 10373 26624 10437 26628
rect 10453 26684 10517 26688
rect 10453 26628 10457 26684
rect 10457 26628 10513 26684
rect 10513 26628 10517 26684
rect 10453 26624 10517 26628
rect 19474 26684 19538 26688
rect 19474 26628 19478 26684
rect 19478 26628 19534 26684
rect 19534 26628 19538 26684
rect 19474 26624 19538 26628
rect 19554 26684 19618 26688
rect 19554 26628 19558 26684
rect 19558 26628 19614 26684
rect 19614 26628 19618 26684
rect 19554 26624 19618 26628
rect 19634 26684 19698 26688
rect 19634 26628 19638 26684
rect 19638 26628 19694 26684
rect 19694 26628 19698 26684
rect 19634 26624 19698 26628
rect 19714 26684 19778 26688
rect 19714 26628 19718 26684
rect 19718 26628 19774 26684
rect 19774 26628 19778 26684
rect 19714 26624 19778 26628
rect 5582 26140 5646 26144
rect 5582 26084 5586 26140
rect 5586 26084 5642 26140
rect 5642 26084 5646 26140
rect 5582 26080 5646 26084
rect 5662 26140 5726 26144
rect 5662 26084 5666 26140
rect 5666 26084 5722 26140
rect 5722 26084 5726 26140
rect 5662 26080 5726 26084
rect 5742 26140 5806 26144
rect 5742 26084 5746 26140
rect 5746 26084 5802 26140
rect 5802 26084 5806 26140
rect 5742 26080 5806 26084
rect 5822 26140 5886 26144
rect 5822 26084 5826 26140
rect 5826 26084 5882 26140
rect 5882 26084 5886 26140
rect 5822 26080 5886 26084
rect 14844 26140 14908 26144
rect 14844 26084 14848 26140
rect 14848 26084 14904 26140
rect 14904 26084 14908 26140
rect 14844 26080 14908 26084
rect 14924 26140 14988 26144
rect 14924 26084 14928 26140
rect 14928 26084 14984 26140
rect 14984 26084 14988 26140
rect 14924 26080 14988 26084
rect 15004 26140 15068 26144
rect 15004 26084 15008 26140
rect 15008 26084 15064 26140
rect 15064 26084 15068 26140
rect 15004 26080 15068 26084
rect 15084 26140 15148 26144
rect 15084 26084 15088 26140
rect 15088 26084 15144 26140
rect 15144 26084 15148 26140
rect 15084 26080 15148 26084
rect 24105 26140 24169 26144
rect 24105 26084 24109 26140
rect 24109 26084 24165 26140
rect 24165 26084 24169 26140
rect 24105 26080 24169 26084
rect 24185 26140 24249 26144
rect 24185 26084 24189 26140
rect 24189 26084 24245 26140
rect 24245 26084 24249 26140
rect 24185 26080 24249 26084
rect 24265 26140 24329 26144
rect 24265 26084 24269 26140
rect 24269 26084 24325 26140
rect 24325 26084 24329 26140
rect 24265 26080 24329 26084
rect 24345 26140 24409 26144
rect 24345 26084 24349 26140
rect 24349 26084 24405 26140
rect 24405 26084 24409 26140
rect 24345 26080 24409 26084
rect 10213 25596 10277 25600
rect 10213 25540 10217 25596
rect 10217 25540 10273 25596
rect 10273 25540 10277 25596
rect 10213 25536 10277 25540
rect 10293 25596 10357 25600
rect 10293 25540 10297 25596
rect 10297 25540 10353 25596
rect 10353 25540 10357 25596
rect 10293 25536 10357 25540
rect 10373 25596 10437 25600
rect 10373 25540 10377 25596
rect 10377 25540 10433 25596
rect 10433 25540 10437 25596
rect 10373 25536 10437 25540
rect 10453 25596 10517 25600
rect 10453 25540 10457 25596
rect 10457 25540 10513 25596
rect 10513 25540 10517 25596
rect 10453 25536 10517 25540
rect 19474 25596 19538 25600
rect 19474 25540 19478 25596
rect 19478 25540 19534 25596
rect 19534 25540 19538 25596
rect 19474 25536 19538 25540
rect 19554 25596 19618 25600
rect 19554 25540 19558 25596
rect 19558 25540 19614 25596
rect 19614 25540 19618 25596
rect 19554 25536 19618 25540
rect 19634 25596 19698 25600
rect 19634 25540 19638 25596
rect 19638 25540 19694 25596
rect 19694 25540 19698 25596
rect 19634 25536 19698 25540
rect 19714 25596 19778 25600
rect 19714 25540 19718 25596
rect 19718 25540 19774 25596
rect 19774 25540 19778 25596
rect 19714 25536 19778 25540
rect 5582 25052 5646 25056
rect 5582 24996 5586 25052
rect 5586 24996 5642 25052
rect 5642 24996 5646 25052
rect 5582 24992 5646 24996
rect 5662 25052 5726 25056
rect 5662 24996 5666 25052
rect 5666 24996 5722 25052
rect 5722 24996 5726 25052
rect 5662 24992 5726 24996
rect 5742 25052 5806 25056
rect 5742 24996 5746 25052
rect 5746 24996 5802 25052
rect 5802 24996 5806 25052
rect 5742 24992 5806 24996
rect 5822 25052 5886 25056
rect 5822 24996 5826 25052
rect 5826 24996 5882 25052
rect 5882 24996 5886 25052
rect 5822 24992 5886 24996
rect 14844 25052 14908 25056
rect 14844 24996 14848 25052
rect 14848 24996 14904 25052
rect 14904 24996 14908 25052
rect 14844 24992 14908 24996
rect 14924 25052 14988 25056
rect 14924 24996 14928 25052
rect 14928 24996 14984 25052
rect 14984 24996 14988 25052
rect 14924 24992 14988 24996
rect 15004 25052 15068 25056
rect 15004 24996 15008 25052
rect 15008 24996 15064 25052
rect 15064 24996 15068 25052
rect 15004 24992 15068 24996
rect 15084 25052 15148 25056
rect 15084 24996 15088 25052
rect 15088 24996 15144 25052
rect 15144 24996 15148 25052
rect 15084 24992 15148 24996
rect 24105 25052 24169 25056
rect 24105 24996 24109 25052
rect 24109 24996 24165 25052
rect 24165 24996 24169 25052
rect 24105 24992 24169 24996
rect 24185 25052 24249 25056
rect 24185 24996 24189 25052
rect 24189 24996 24245 25052
rect 24245 24996 24249 25052
rect 24185 24992 24249 24996
rect 24265 25052 24329 25056
rect 24265 24996 24269 25052
rect 24269 24996 24325 25052
rect 24325 24996 24329 25052
rect 24265 24992 24329 24996
rect 24345 25052 24409 25056
rect 24345 24996 24349 25052
rect 24349 24996 24405 25052
rect 24405 24996 24409 25052
rect 24345 24992 24409 24996
rect 10213 24508 10277 24512
rect 10213 24452 10217 24508
rect 10217 24452 10273 24508
rect 10273 24452 10277 24508
rect 10213 24448 10277 24452
rect 10293 24508 10357 24512
rect 10293 24452 10297 24508
rect 10297 24452 10353 24508
rect 10353 24452 10357 24508
rect 10293 24448 10357 24452
rect 10373 24508 10437 24512
rect 10373 24452 10377 24508
rect 10377 24452 10433 24508
rect 10433 24452 10437 24508
rect 10373 24448 10437 24452
rect 10453 24508 10517 24512
rect 10453 24452 10457 24508
rect 10457 24452 10513 24508
rect 10513 24452 10517 24508
rect 10453 24448 10517 24452
rect 19474 24508 19538 24512
rect 19474 24452 19478 24508
rect 19478 24452 19534 24508
rect 19534 24452 19538 24508
rect 19474 24448 19538 24452
rect 19554 24508 19618 24512
rect 19554 24452 19558 24508
rect 19558 24452 19614 24508
rect 19614 24452 19618 24508
rect 19554 24448 19618 24452
rect 19634 24508 19698 24512
rect 19634 24452 19638 24508
rect 19638 24452 19694 24508
rect 19694 24452 19698 24508
rect 19634 24448 19698 24452
rect 19714 24508 19778 24512
rect 19714 24452 19718 24508
rect 19718 24452 19774 24508
rect 19774 24452 19778 24508
rect 19714 24448 19778 24452
rect 5582 23964 5646 23968
rect 5582 23908 5586 23964
rect 5586 23908 5642 23964
rect 5642 23908 5646 23964
rect 5582 23904 5646 23908
rect 5662 23964 5726 23968
rect 5662 23908 5666 23964
rect 5666 23908 5722 23964
rect 5722 23908 5726 23964
rect 5662 23904 5726 23908
rect 5742 23964 5806 23968
rect 5742 23908 5746 23964
rect 5746 23908 5802 23964
rect 5802 23908 5806 23964
rect 5742 23904 5806 23908
rect 5822 23964 5886 23968
rect 5822 23908 5826 23964
rect 5826 23908 5882 23964
rect 5882 23908 5886 23964
rect 5822 23904 5886 23908
rect 14844 23964 14908 23968
rect 14844 23908 14848 23964
rect 14848 23908 14904 23964
rect 14904 23908 14908 23964
rect 14844 23904 14908 23908
rect 14924 23964 14988 23968
rect 14924 23908 14928 23964
rect 14928 23908 14984 23964
rect 14984 23908 14988 23964
rect 14924 23904 14988 23908
rect 15004 23964 15068 23968
rect 15004 23908 15008 23964
rect 15008 23908 15064 23964
rect 15064 23908 15068 23964
rect 15004 23904 15068 23908
rect 15084 23964 15148 23968
rect 15084 23908 15088 23964
rect 15088 23908 15144 23964
rect 15144 23908 15148 23964
rect 15084 23904 15148 23908
rect 24105 23964 24169 23968
rect 24105 23908 24109 23964
rect 24109 23908 24165 23964
rect 24165 23908 24169 23964
rect 24105 23904 24169 23908
rect 24185 23964 24249 23968
rect 24185 23908 24189 23964
rect 24189 23908 24245 23964
rect 24245 23908 24249 23964
rect 24185 23904 24249 23908
rect 24265 23964 24329 23968
rect 24265 23908 24269 23964
rect 24269 23908 24325 23964
rect 24325 23908 24329 23964
rect 24265 23904 24329 23908
rect 24345 23964 24409 23968
rect 24345 23908 24349 23964
rect 24349 23908 24405 23964
rect 24405 23908 24409 23964
rect 24345 23904 24409 23908
rect 10213 23420 10277 23424
rect 10213 23364 10217 23420
rect 10217 23364 10273 23420
rect 10273 23364 10277 23420
rect 10213 23360 10277 23364
rect 10293 23420 10357 23424
rect 10293 23364 10297 23420
rect 10297 23364 10353 23420
rect 10353 23364 10357 23420
rect 10293 23360 10357 23364
rect 10373 23420 10437 23424
rect 10373 23364 10377 23420
rect 10377 23364 10433 23420
rect 10433 23364 10437 23420
rect 10373 23360 10437 23364
rect 10453 23420 10517 23424
rect 10453 23364 10457 23420
rect 10457 23364 10513 23420
rect 10513 23364 10517 23420
rect 10453 23360 10517 23364
rect 19474 23420 19538 23424
rect 19474 23364 19478 23420
rect 19478 23364 19534 23420
rect 19534 23364 19538 23420
rect 19474 23360 19538 23364
rect 19554 23420 19618 23424
rect 19554 23364 19558 23420
rect 19558 23364 19614 23420
rect 19614 23364 19618 23420
rect 19554 23360 19618 23364
rect 19634 23420 19698 23424
rect 19634 23364 19638 23420
rect 19638 23364 19694 23420
rect 19694 23364 19698 23420
rect 19634 23360 19698 23364
rect 19714 23420 19778 23424
rect 19714 23364 19718 23420
rect 19718 23364 19774 23420
rect 19774 23364 19778 23420
rect 19714 23360 19778 23364
rect 5582 22876 5646 22880
rect 5582 22820 5586 22876
rect 5586 22820 5642 22876
rect 5642 22820 5646 22876
rect 5582 22816 5646 22820
rect 5662 22876 5726 22880
rect 5662 22820 5666 22876
rect 5666 22820 5722 22876
rect 5722 22820 5726 22876
rect 5662 22816 5726 22820
rect 5742 22876 5806 22880
rect 5742 22820 5746 22876
rect 5746 22820 5802 22876
rect 5802 22820 5806 22876
rect 5742 22816 5806 22820
rect 5822 22876 5886 22880
rect 5822 22820 5826 22876
rect 5826 22820 5882 22876
rect 5882 22820 5886 22876
rect 5822 22816 5886 22820
rect 14844 22876 14908 22880
rect 14844 22820 14848 22876
rect 14848 22820 14904 22876
rect 14904 22820 14908 22876
rect 14844 22816 14908 22820
rect 14924 22876 14988 22880
rect 14924 22820 14928 22876
rect 14928 22820 14984 22876
rect 14984 22820 14988 22876
rect 14924 22816 14988 22820
rect 15004 22876 15068 22880
rect 15004 22820 15008 22876
rect 15008 22820 15064 22876
rect 15064 22820 15068 22876
rect 15004 22816 15068 22820
rect 15084 22876 15148 22880
rect 15084 22820 15088 22876
rect 15088 22820 15144 22876
rect 15144 22820 15148 22876
rect 15084 22816 15148 22820
rect 24105 22876 24169 22880
rect 24105 22820 24109 22876
rect 24109 22820 24165 22876
rect 24165 22820 24169 22876
rect 24105 22816 24169 22820
rect 24185 22876 24249 22880
rect 24185 22820 24189 22876
rect 24189 22820 24245 22876
rect 24245 22820 24249 22876
rect 24185 22816 24249 22820
rect 24265 22876 24329 22880
rect 24265 22820 24269 22876
rect 24269 22820 24325 22876
rect 24325 22820 24329 22876
rect 24265 22816 24329 22820
rect 24345 22876 24409 22880
rect 24345 22820 24349 22876
rect 24349 22820 24405 22876
rect 24405 22820 24409 22876
rect 24345 22816 24409 22820
rect 10213 22332 10277 22336
rect 10213 22276 10217 22332
rect 10217 22276 10273 22332
rect 10273 22276 10277 22332
rect 10213 22272 10277 22276
rect 10293 22332 10357 22336
rect 10293 22276 10297 22332
rect 10297 22276 10353 22332
rect 10353 22276 10357 22332
rect 10293 22272 10357 22276
rect 10373 22332 10437 22336
rect 10373 22276 10377 22332
rect 10377 22276 10433 22332
rect 10433 22276 10437 22332
rect 10373 22272 10437 22276
rect 10453 22332 10517 22336
rect 10453 22276 10457 22332
rect 10457 22276 10513 22332
rect 10513 22276 10517 22332
rect 10453 22272 10517 22276
rect 19474 22332 19538 22336
rect 19474 22276 19478 22332
rect 19478 22276 19534 22332
rect 19534 22276 19538 22332
rect 19474 22272 19538 22276
rect 19554 22332 19618 22336
rect 19554 22276 19558 22332
rect 19558 22276 19614 22332
rect 19614 22276 19618 22332
rect 19554 22272 19618 22276
rect 19634 22332 19698 22336
rect 19634 22276 19638 22332
rect 19638 22276 19694 22332
rect 19694 22276 19698 22332
rect 19634 22272 19698 22276
rect 19714 22332 19778 22336
rect 19714 22276 19718 22332
rect 19718 22276 19774 22332
rect 19774 22276 19778 22332
rect 19714 22272 19778 22276
rect 5582 21788 5646 21792
rect 5582 21732 5586 21788
rect 5586 21732 5642 21788
rect 5642 21732 5646 21788
rect 5582 21728 5646 21732
rect 5662 21788 5726 21792
rect 5662 21732 5666 21788
rect 5666 21732 5722 21788
rect 5722 21732 5726 21788
rect 5662 21728 5726 21732
rect 5742 21788 5806 21792
rect 5742 21732 5746 21788
rect 5746 21732 5802 21788
rect 5802 21732 5806 21788
rect 5742 21728 5806 21732
rect 5822 21788 5886 21792
rect 5822 21732 5826 21788
rect 5826 21732 5882 21788
rect 5882 21732 5886 21788
rect 5822 21728 5886 21732
rect 14844 21788 14908 21792
rect 14844 21732 14848 21788
rect 14848 21732 14904 21788
rect 14904 21732 14908 21788
rect 14844 21728 14908 21732
rect 14924 21788 14988 21792
rect 14924 21732 14928 21788
rect 14928 21732 14984 21788
rect 14984 21732 14988 21788
rect 14924 21728 14988 21732
rect 15004 21788 15068 21792
rect 15004 21732 15008 21788
rect 15008 21732 15064 21788
rect 15064 21732 15068 21788
rect 15004 21728 15068 21732
rect 15084 21788 15148 21792
rect 15084 21732 15088 21788
rect 15088 21732 15144 21788
rect 15144 21732 15148 21788
rect 15084 21728 15148 21732
rect 24105 21788 24169 21792
rect 24105 21732 24109 21788
rect 24109 21732 24165 21788
rect 24165 21732 24169 21788
rect 24105 21728 24169 21732
rect 24185 21788 24249 21792
rect 24185 21732 24189 21788
rect 24189 21732 24245 21788
rect 24245 21732 24249 21788
rect 24185 21728 24249 21732
rect 24265 21788 24329 21792
rect 24265 21732 24269 21788
rect 24269 21732 24325 21788
rect 24325 21732 24329 21788
rect 24265 21728 24329 21732
rect 24345 21788 24409 21792
rect 24345 21732 24349 21788
rect 24349 21732 24405 21788
rect 24405 21732 24409 21788
rect 24345 21728 24409 21732
rect 10213 21244 10277 21248
rect 10213 21188 10217 21244
rect 10217 21188 10273 21244
rect 10273 21188 10277 21244
rect 10213 21184 10277 21188
rect 10293 21244 10357 21248
rect 10293 21188 10297 21244
rect 10297 21188 10353 21244
rect 10353 21188 10357 21244
rect 10293 21184 10357 21188
rect 10373 21244 10437 21248
rect 10373 21188 10377 21244
rect 10377 21188 10433 21244
rect 10433 21188 10437 21244
rect 10373 21184 10437 21188
rect 10453 21244 10517 21248
rect 10453 21188 10457 21244
rect 10457 21188 10513 21244
rect 10513 21188 10517 21244
rect 10453 21184 10517 21188
rect 19474 21244 19538 21248
rect 19474 21188 19478 21244
rect 19478 21188 19534 21244
rect 19534 21188 19538 21244
rect 19474 21184 19538 21188
rect 19554 21244 19618 21248
rect 19554 21188 19558 21244
rect 19558 21188 19614 21244
rect 19614 21188 19618 21244
rect 19554 21184 19618 21188
rect 19634 21244 19698 21248
rect 19634 21188 19638 21244
rect 19638 21188 19694 21244
rect 19694 21188 19698 21244
rect 19634 21184 19698 21188
rect 19714 21244 19778 21248
rect 19714 21188 19718 21244
rect 19718 21188 19774 21244
rect 19774 21188 19778 21244
rect 19714 21184 19778 21188
rect 5582 20700 5646 20704
rect 5582 20644 5586 20700
rect 5586 20644 5642 20700
rect 5642 20644 5646 20700
rect 5582 20640 5646 20644
rect 5662 20700 5726 20704
rect 5662 20644 5666 20700
rect 5666 20644 5722 20700
rect 5722 20644 5726 20700
rect 5662 20640 5726 20644
rect 5742 20700 5806 20704
rect 5742 20644 5746 20700
rect 5746 20644 5802 20700
rect 5802 20644 5806 20700
rect 5742 20640 5806 20644
rect 5822 20700 5886 20704
rect 5822 20644 5826 20700
rect 5826 20644 5882 20700
rect 5882 20644 5886 20700
rect 5822 20640 5886 20644
rect 14844 20700 14908 20704
rect 14844 20644 14848 20700
rect 14848 20644 14904 20700
rect 14904 20644 14908 20700
rect 14844 20640 14908 20644
rect 14924 20700 14988 20704
rect 14924 20644 14928 20700
rect 14928 20644 14984 20700
rect 14984 20644 14988 20700
rect 14924 20640 14988 20644
rect 15004 20700 15068 20704
rect 15004 20644 15008 20700
rect 15008 20644 15064 20700
rect 15064 20644 15068 20700
rect 15004 20640 15068 20644
rect 15084 20700 15148 20704
rect 15084 20644 15088 20700
rect 15088 20644 15144 20700
rect 15144 20644 15148 20700
rect 15084 20640 15148 20644
rect 24105 20700 24169 20704
rect 24105 20644 24109 20700
rect 24109 20644 24165 20700
rect 24165 20644 24169 20700
rect 24105 20640 24169 20644
rect 24185 20700 24249 20704
rect 24185 20644 24189 20700
rect 24189 20644 24245 20700
rect 24245 20644 24249 20700
rect 24185 20640 24249 20644
rect 24265 20700 24329 20704
rect 24265 20644 24269 20700
rect 24269 20644 24325 20700
rect 24325 20644 24329 20700
rect 24265 20640 24329 20644
rect 24345 20700 24409 20704
rect 24345 20644 24349 20700
rect 24349 20644 24405 20700
rect 24405 20644 24409 20700
rect 24345 20640 24409 20644
rect 10213 20156 10277 20160
rect 10213 20100 10217 20156
rect 10217 20100 10273 20156
rect 10273 20100 10277 20156
rect 10213 20096 10277 20100
rect 10293 20156 10357 20160
rect 10293 20100 10297 20156
rect 10297 20100 10353 20156
rect 10353 20100 10357 20156
rect 10293 20096 10357 20100
rect 10373 20156 10437 20160
rect 10373 20100 10377 20156
rect 10377 20100 10433 20156
rect 10433 20100 10437 20156
rect 10373 20096 10437 20100
rect 10453 20156 10517 20160
rect 10453 20100 10457 20156
rect 10457 20100 10513 20156
rect 10513 20100 10517 20156
rect 10453 20096 10517 20100
rect 19474 20156 19538 20160
rect 19474 20100 19478 20156
rect 19478 20100 19534 20156
rect 19534 20100 19538 20156
rect 19474 20096 19538 20100
rect 19554 20156 19618 20160
rect 19554 20100 19558 20156
rect 19558 20100 19614 20156
rect 19614 20100 19618 20156
rect 19554 20096 19618 20100
rect 19634 20156 19698 20160
rect 19634 20100 19638 20156
rect 19638 20100 19694 20156
rect 19694 20100 19698 20156
rect 19634 20096 19698 20100
rect 19714 20156 19778 20160
rect 19714 20100 19718 20156
rect 19718 20100 19774 20156
rect 19774 20100 19778 20156
rect 19714 20096 19778 20100
rect 5582 19612 5646 19616
rect 5582 19556 5586 19612
rect 5586 19556 5642 19612
rect 5642 19556 5646 19612
rect 5582 19552 5646 19556
rect 5662 19612 5726 19616
rect 5662 19556 5666 19612
rect 5666 19556 5722 19612
rect 5722 19556 5726 19612
rect 5662 19552 5726 19556
rect 5742 19612 5806 19616
rect 5742 19556 5746 19612
rect 5746 19556 5802 19612
rect 5802 19556 5806 19612
rect 5742 19552 5806 19556
rect 5822 19612 5886 19616
rect 5822 19556 5826 19612
rect 5826 19556 5882 19612
rect 5882 19556 5886 19612
rect 5822 19552 5886 19556
rect 14844 19612 14908 19616
rect 14844 19556 14848 19612
rect 14848 19556 14904 19612
rect 14904 19556 14908 19612
rect 14844 19552 14908 19556
rect 14924 19612 14988 19616
rect 14924 19556 14928 19612
rect 14928 19556 14984 19612
rect 14984 19556 14988 19612
rect 14924 19552 14988 19556
rect 15004 19612 15068 19616
rect 15004 19556 15008 19612
rect 15008 19556 15064 19612
rect 15064 19556 15068 19612
rect 15004 19552 15068 19556
rect 15084 19612 15148 19616
rect 15084 19556 15088 19612
rect 15088 19556 15144 19612
rect 15144 19556 15148 19612
rect 15084 19552 15148 19556
rect 24105 19612 24169 19616
rect 24105 19556 24109 19612
rect 24109 19556 24165 19612
rect 24165 19556 24169 19612
rect 24105 19552 24169 19556
rect 24185 19612 24249 19616
rect 24185 19556 24189 19612
rect 24189 19556 24245 19612
rect 24245 19556 24249 19612
rect 24185 19552 24249 19556
rect 24265 19612 24329 19616
rect 24265 19556 24269 19612
rect 24269 19556 24325 19612
rect 24325 19556 24329 19612
rect 24265 19552 24329 19556
rect 24345 19612 24409 19616
rect 24345 19556 24349 19612
rect 24349 19556 24405 19612
rect 24405 19556 24409 19612
rect 24345 19552 24409 19556
rect 10213 19068 10277 19072
rect 10213 19012 10217 19068
rect 10217 19012 10273 19068
rect 10273 19012 10277 19068
rect 10213 19008 10277 19012
rect 10293 19068 10357 19072
rect 10293 19012 10297 19068
rect 10297 19012 10353 19068
rect 10353 19012 10357 19068
rect 10293 19008 10357 19012
rect 10373 19068 10437 19072
rect 10373 19012 10377 19068
rect 10377 19012 10433 19068
rect 10433 19012 10437 19068
rect 10373 19008 10437 19012
rect 10453 19068 10517 19072
rect 10453 19012 10457 19068
rect 10457 19012 10513 19068
rect 10513 19012 10517 19068
rect 10453 19008 10517 19012
rect 19474 19068 19538 19072
rect 19474 19012 19478 19068
rect 19478 19012 19534 19068
rect 19534 19012 19538 19068
rect 19474 19008 19538 19012
rect 19554 19068 19618 19072
rect 19554 19012 19558 19068
rect 19558 19012 19614 19068
rect 19614 19012 19618 19068
rect 19554 19008 19618 19012
rect 19634 19068 19698 19072
rect 19634 19012 19638 19068
rect 19638 19012 19694 19068
rect 19694 19012 19698 19068
rect 19634 19008 19698 19012
rect 19714 19068 19778 19072
rect 19714 19012 19718 19068
rect 19718 19012 19774 19068
rect 19774 19012 19778 19068
rect 19714 19008 19778 19012
rect 5582 18524 5646 18528
rect 5582 18468 5586 18524
rect 5586 18468 5642 18524
rect 5642 18468 5646 18524
rect 5582 18464 5646 18468
rect 5662 18524 5726 18528
rect 5662 18468 5666 18524
rect 5666 18468 5722 18524
rect 5722 18468 5726 18524
rect 5662 18464 5726 18468
rect 5742 18524 5806 18528
rect 5742 18468 5746 18524
rect 5746 18468 5802 18524
rect 5802 18468 5806 18524
rect 5742 18464 5806 18468
rect 5822 18524 5886 18528
rect 5822 18468 5826 18524
rect 5826 18468 5882 18524
rect 5882 18468 5886 18524
rect 5822 18464 5886 18468
rect 14844 18524 14908 18528
rect 14844 18468 14848 18524
rect 14848 18468 14904 18524
rect 14904 18468 14908 18524
rect 14844 18464 14908 18468
rect 14924 18524 14988 18528
rect 14924 18468 14928 18524
rect 14928 18468 14984 18524
rect 14984 18468 14988 18524
rect 14924 18464 14988 18468
rect 15004 18524 15068 18528
rect 15004 18468 15008 18524
rect 15008 18468 15064 18524
rect 15064 18468 15068 18524
rect 15004 18464 15068 18468
rect 15084 18524 15148 18528
rect 15084 18468 15088 18524
rect 15088 18468 15144 18524
rect 15144 18468 15148 18524
rect 15084 18464 15148 18468
rect 24105 18524 24169 18528
rect 24105 18468 24109 18524
rect 24109 18468 24165 18524
rect 24165 18468 24169 18524
rect 24105 18464 24169 18468
rect 24185 18524 24249 18528
rect 24185 18468 24189 18524
rect 24189 18468 24245 18524
rect 24245 18468 24249 18524
rect 24185 18464 24249 18468
rect 24265 18524 24329 18528
rect 24265 18468 24269 18524
rect 24269 18468 24325 18524
rect 24325 18468 24329 18524
rect 24265 18464 24329 18468
rect 24345 18524 24409 18528
rect 24345 18468 24349 18524
rect 24349 18468 24405 18524
rect 24405 18468 24409 18524
rect 24345 18464 24409 18468
rect 10213 17980 10277 17984
rect 10213 17924 10217 17980
rect 10217 17924 10273 17980
rect 10273 17924 10277 17980
rect 10213 17920 10277 17924
rect 10293 17980 10357 17984
rect 10293 17924 10297 17980
rect 10297 17924 10353 17980
rect 10353 17924 10357 17980
rect 10293 17920 10357 17924
rect 10373 17980 10437 17984
rect 10373 17924 10377 17980
rect 10377 17924 10433 17980
rect 10433 17924 10437 17980
rect 10373 17920 10437 17924
rect 10453 17980 10517 17984
rect 10453 17924 10457 17980
rect 10457 17924 10513 17980
rect 10513 17924 10517 17980
rect 10453 17920 10517 17924
rect 19474 17980 19538 17984
rect 19474 17924 19478 17980
rect 19478 17924 19534 17980
rect 19534 17924 19538 17980
rect 19474 17920 19538 17924
rect 19554 17980 19618 17984
rect 19554 17924 19558 17980
rect 19558 17924 19614 17980
rect 19614 17924 19618 17980
rect 19554 17920 19618 17924
rect 19634 17980 19698 17984
rect 19634 17924 19638 17980
rect 19638 17924 19694 17980
rect 19694 17924 19698 17980
rect 19634 17920 19698 17924
rect 19714 17980 19778 17984
rect 19714 17924 19718 17980
rect 19718 17924 19774 17980
rect 19774 17924 19778 17980
rect 19714 17920 19778 17924
rect 5582 17436 5646 17440
rect 5582 17380 5586 17436
rect 5586 17380 5642 17436
rect 5642 17380 5646 17436
rect 5582 17376 5646 17380
rect 5662 17436 5726 17440
rect 5662 17380 5666 17436
rect 5666 17380 5722 17436
rect 5722 17380 5726 17436
rect 5662 17376 5726 17380
rect 5742 17436 5806 17440
rect 5742 17380 5746 17436
rect 5746 17380 5802 17436
rect 5802 17380 5806 17436
rect 5742 17376 5806 17380
rect 5822 17436 5886 17440
rect 5822 17380 5826 17436
rect 5826 17380 5882 17436
rect 5882 17380 5886 17436
rect 5822 17376 5886 17380
rect 14844 17436 14908 17440
rect 14844 17380 14848 17436
rect 14848 17380 14904 17436
rect 14904 17380 14908 17436
rect 14844 17376 14908 17380
rect 14924 17436 14988 17440
rect 14924 17380 14928 17436
rect 14928 17380 14984 17436
rect 14984 17380 14988 17436
rect 14924 17376 14988 17380
rect 15004 17436 15068 17440
rect 15004 17380 15008 17436
rect 15008 17380 15064 17436
rect 15064 17380 15068 17436
rect 15004 17376 15068 17380
rect 15084 17436 15148 17440
rect 15084 17380 15088 17436
rect 15088 17380 15144 17436
rect 15144 17380 15148 17436
rect 15084 17376 15148 17380
rect 24105 17436 24169 17440
rect 24105 17380 24109 17436
rect 24109 17380 24165 17436
rect 24165 17380 24169 17436
rect 24105 17376 24169 17380
rect 24185 17436 24249 17440
rect 24185 17380 24189 17436
rect 24189 17380 24245 17436
rect 24245 17380 24249 17436
rect 24185 17376 24249 17380
rect 24265 17436 24329 17440
rect 24265 17380 24269 17436
rect 24269 17380 24325 17436
rect 24325 17380 24329 17436
rect 24265 17376 24329 17380
rect 24345 17436 24409 17440
rect 24345 17380 24349 17436
rect 24349 17380 24405 17436
rect 24405 17380 24409 17436
rect 24345 17376 24409 17380
rect 10213 16892 10277 16896
rect 10213 16836 10217 16892
rect 10217 16836 10273 16892
rect 10273 16836 10277 16892
rect 10213 16832 10277 16836
rect 10293 16892 10357 16896
rect 10293 16836 10297 16892
rect 10297 16836 10353 16892
rect 10353 16836 10357 16892
rect 10293 16832 10357 16836
rect 10373 16892 10437 16896
rect 10373 16836 10377 16892
rect 10377 16836 10433 16892
rect 10433 16836 10437 16892
rect 10373 16832 10437 16836
rect 10453 16892 10517 16896
rect 10453 16836 10457 16892
rect 10457 16836 10513 16892
rect 10513 16836 10517 16892
rect 10453 16832 10517 16836
rect 19474 16892 19538 16896
rect 19474 16836 19478 16892
rect 19478 16836 19534 16892
rect 19534 16836 19538 16892
rect 19474 16832 19538 16836
rect 19554 16892 19618 16896
rect 19554 16836 19558 16892
rect 19558 16836 19614 16892
rect 19614 16836 19618 16892
rect 19554 16832 19618 16836
rect 19634 16892 19698 16896
rect 19634 16836 19638 16892
rect 19638 16836 19694 16892
rect 19694 16836 19698 16892
rect 19634 16832 19698 16836
rect 19714 16892 19778 16896
rect 19714 16836 19718 16892
rect 19718 16836 19774 16892
rect 19774 16836 19778 16892
rect 19714 16832 19778 16836
rect 5582 16348 5646 16352
rect 5582 16292 5586 16348
rect 5586 16292 5642 16348
rect 5642 16292 5646 16348
rect 5582 16288 5646 16292
rect 5662 16348 5726 16352
rect 5662 16292 5666 16348
rect 5666 16292 5722 16348
rect 5722 16292 5726 16348
rect 5662 16288 5726 16292
rect 5742 16348 5806 16352
rect 5742 16292 5746 16348
rect 5746 16292 5802 16348
rect 5802 16292 5806 16348
rect 5742 16288 5806 16292
rect 5822 16348 5886 16352
rect 5822 16292 5826 16348
rect 5826 16292 5882 16348
rect 5882 16292 5886 16348
rect 5822 16288 5886 16292
rect 14844 16348 14908 16352
rect 14844 16292 14848 16348
rect 14848 16292 14904 16348
rect 14904 16292 14908 16348
rect 14844 16288 14908 16292
rect 14924 16348 14988 16352
rect 14924 16292 14928 16348
rect 14928 16292 14984 16348
rect 14984 16292 14988 16348
rect 14924 16288 14988 16292
rect 15004 16348 15068 16352
rect 15004 16292 15008 16348
rect 15008 16292 15064 16348
rect 15064 16292 15068 16348
rect 15004 16288 15068 16292
rect 15084 16348 15148 16352
rect 15084 16292 15088 16348
rect 15088 16292 15144 16348
rect 15144 16292 15148 16348
rect 15084 16288 15148 16292
rect 24105 16348 24169 16352
rect 24105 16292 24109 16348
rect 24109 16292 24165 16348
rect 24165 16292 24169 16348
rect 24105 16288 24169 16292
rect 24185 16348 24249 16352
rect 24185 16292 24189 16348
rect 24189 16292 24245 16348
rect 24245 16292 24249 16348
rect 24185 16288 24249 16292
rect 24265 16348 24329 16352
rect 24265 16292 24269 16348
rect 24269 16292 24325 16348
rect 24325 16292 24329 16348
rect 24265 16288 24329 16292
rect 24345 16348 24409 16352
rect 24345 16292 24349 16348
rect 24349 16292 24405 16348
rect 24405 16292 24409 16348
rect 24345 16288 24409 16292
rect 10213 15804 10277 15808
rect 10213 15748 10217 15804
rect 10217 15748 10273 15804
rect 10273 15748 10277 15804
rect 10213 15744 10277 15748
rect 10293 15804 10357 15808
rect 10293 15748 10297 15804
rect 10297 15748 10353 15804
rect 10353 15748 10357 15804
rect 10293 15744 10357 15748
rect 10373 15804 10437 15808
rect 10373 15748 10377 15804
rect 10377 15748 10433 15804
rect 10433 15748 10437 15804
rect 10373 15744 10437 15748
rect 10453 15804 10517 15808
rect 10453 15748 10457 15804
rect 10457 15748 10513 15804
rect 10513 15748 10517 15804
rect 10453 15744 10517 15748
rect 19474 15804 19538 15808
rect 19474 15748 19478 15804
rect 19478 15748 19534 15804
rect 19534 15748 19538 15804
rect 19474 15744 19538 15748
rect 19554 15804 19618 15808
rect 19554 15748 19558 15804
rect 19558 15748 19614 15804
rect 19614 15748 19618 15804
rect 19554 15744 19618 15748
rect 19634 15804 19698 15808
rect 19634 15748 19638 15804
rect 19638 15748 19694 15804
rect 19694 15748 19698 15804
rect 19634 15744 19698 15748
rect 19714 15804 19778 15808
rect 19714 15748 19718 15804
rect 19718 15748 19774 15804
rect 19774 15748 19778 15804
rect 19714 15744 19778 15748
rect 5582 15260 5646 15264
rect 5582 15204 5586 15260
rect 5586 15204 5642 15260
rect 5642 15204 5646 15260
rect 5582 15200 5646 15204
rect 5662 15260 5726 15264
rect 5662 15204 5666 15260
rect 5666 15204 5722 15260
rect 5722 15204 5726 15260
rect 5662 15200 5726 15204
rect 5742 15260 5806 15264
rect 5742 15204 5746 15260
rect 5746 15204 5802 15260
rect 5802 15204 5806 15260
rect 5742 15200 5806 15204
rect 5822 15260 5886 15264
rect 5822 15204 5826 15260
rect 5826 15204 5882 15260
rect 5882 15204 5886 15260
rect 5822 15200 5886 15204
rect 14844 15260 14908 15264
rect 14844 15204 14848 15260
rect 14848 15204 14904 15260
rect 14904 15204 14908 15260
rect 14844 15200 14908 15204
rect 14924 15260 14988 15264
rect 14924 15204 14928 15260
rect 14928 15204 14984 15260
rect 14984 15204 14988 15260
rect 14924 15200 14988 15204
rect 15004 15260 15068 15264
rect 15004 15204 15008 15260
rect 15008 15204 15064 15260
rect 15064 15204 15068 15260
rect 15004 15200 15068 15204
rect 15084 15260 15148 15264
rect 15084 15204 15088 15260
rect 15088 15204 15144 15260
rect 15144 15204 15148 15260
rect 15084 15200 15148 15204
rect 24105 15260 24169 15264
rect 24105 15204 24109 15260
rect 24109 15204 24165 15260
rect 24165 15204 24169 15260
rect 24105 15200 24169 15204
rect 24185 15260 24249 15264
rect 24185 15204 24189 15260
rect 24189 15204 24245 15260
rect 24245 15204 24249 15260
rect 24185 15200 24249 15204
rect 24265 15260 24329 15264
rect 24265 15204 24269 15260
rect 24269 15204 24325 15260
rect 24325 15204 24329 15260
rect 24265 15200 24329 15204
rect 24345 15260 24409 15264
rect 24345 15204 24349 15260
rect 24349 15204 24405 15260
rect 24405 15204 24409 15260
rect 24345 15200 24409 15204
rect 10213 14716 10277 14720
rect 10213 14660 10217 14716
rect 10217 14660 10273 14716
rect 10273 14660 10277 14716
rect 10213 14656 10277 14660
rect 10293 14716 10357 14720
rect 10293 14660 10297 14716
rect 10297 14660 10353 14716
rect 10353 14660 10357 14716
rect 10293 14656 10357 14660
rect 10373 14716 10437 14720
rect 10373 14660 10377 14716
rect 10377 14660 10433 14716
rect 10433 14660 10437 14716
rect 10373 14656 10437 14660
rect 10453 14716 10517 14720
rect 10453 14660 10457 14716
rect 10457 14660 10513 14716
rect 10513 14660 10517 14716
rect 10453 14656 10517 14660
rect 19474 14716 19538 14720
rect 19474 14660 19478 14716
rect 19478 14660 19534 14716
rect 19534 14660 19538 14716
rect 19474 14656 19538 14660
rect 19554 14716 19618 14720
rect 19554 14660 19558 14716
rect 19558 14660 19614 14716
rect 19614 14660 19618 14716
rect 19554 14656 19618 14660
rect 19634 14716 19698 14720
rect 19634 14660 19638 14716
rect 19638 14660 19694 14716
rect 19694 14660 19698 14716
rect 19634 14656 19698 14660
rect 19714 14716 19778 14720
rect 19714 14660 19718 14716
rect 19718 14660 19774 14716
rect 19774 14660 19778 14716
rect 19714 14656 19778 14660
rect 5582 14172 5646 14176
rect 5582 14116 5586 14172
rect 5586 14116 5642 14172
rect 5642 14116 5646 14172
rect 5582 14112 5646 14116
rect 5662 14172 5726 14176
rect 5662 14116 5666 14172
rect 5666 14116 5722 14172
rect 5722 14116 5726 14172
rect 5662 14112 5726 14116
rect 5742 14172 5806 14176
rect 5742 14116 5746 14172
rect 5746 14116 5802 14172
rect 5802 14116 5806 14172
rect 5742 14112 5806 14116
rect 5822 14172 5886 14176
rect 5822 14116 5826 14172
rect 5826 14116 5882 14172
rect 5882 14116 5886 14172
rect 5822 14112 5886 14116
rect 14844 14172 14908 14176
rect 14844 14116 14848 14172
rect 14848 14116 14904 14172
rect 14904 14116 14908 14172
rect 14844 14112 14908 14116
rect 14924 14172 14988 14176
rect 14924 14116 14928 14172
rect 14928 14116 14984 14172
rect 14984 14116 14988 14172
rect 14924 14112 14988 14116
rect 15004 14172 15068 14176
rect 15004 14116 15008 14172
rect 15008 14116 15064 14172
rect 15064 14116 15068 14172
rect 15004 14112 15068 14116
rect 15084 14172 15148 14176
rect 15084 14116 15088 14172
rect 15088 14116 15144 14172
rect 15144 14116 15148 14172
rect 15084 14112 15148 14116
rect 24105 14172 24169 14176
rect 24105 14116 24109 14172
rect 24109 14116 24165 14172
rect 24165 14116 24169 14172
rect 24105 14112 24169 14116
rect 24185 14172 24249 14176
rect 24185 14116 24189 14172
rect 24189 14116 24245 14172
rect 24245 14116 24249 14172
rect 24185 14112 24249 14116
rect 24265 14172 24329 14176
rect 24265 14116 24269 14172
rect 24269 14116 24325 14172
rect 24325 14116 24329 14172
rect 24265 14112 24329 14116
rect 24345 14172 24409 14176
rect 24345 14116 24349 14172
rect 24349 14116 24405 14172
rect 24405 14116 24409 14172
rect 24345 14112 24409 14116
rect 10213 13628 10277 13632
rect 10213 13572 10217 13628
rect 10217 13572 10273 13628
rect 10273 13572 10277 13628
rect 10213 13568 10277 13572
rect 10293 13628 10357 13632
rect 10293 13572 10297 13628
rect 10297 13572 10353 13628
rect 10353 13572 10357 13628
rect 10293 13568 10357 13572
rect 10373 13628 10437 13632
rect 10373 13572 10377 13628
rect 10377 13572 10433 13628
rect 10433 13572 10437 13628
rect 10373 13568 10437 13572
rect 10453 13628 10517 13632
rect 10453 13572 10457 13628
rect 10457 13572 10513 13628
rect 10513 13572 10517 13628
rect 10453 13568 10517 13572
rect 19474 13628 19538 13632
rect 19474 13572 19478 13628
rect 19478 13572 19534 13628
rect 19534 13572 19538 13628
rect 19474 13568 19538 13572
rect 19554 13628 19618 13632
rect 19554 13572 19558 13628
rect 19558 13572 19614 13628
rect 19614 13572 19618 13628
rect 19554 13568 19618 13572
rect 19634 13628 19698 13632
rect 19634 13572 19638 13628
rect 19638 13572 19694 13628
rect 19694 13572 19698 13628
rect 19634 13568 19698 13572
rect 19714 13628 19778 13632
rect 19714 13572 19718 13628
rect 19718 13572 19774 13628
rect 19774 13572 19778 13628
rect 19714 13568 19778 13572
rect 5582 13084 5646 13088
rect 5582 13028 5586 13084
rect 5586 13028 5642 13084
rect 5642 13028 5646 13084
rect 5582 13024 5646 13028
rect 5662 13084 5726 13088
rect 5662 13028 5666 13084
rect 5666 13028 5722 13084
rect 5722 13028 5726 13084
rect 5662 13024 5726 13028
rect 5742 13084 5806 13088
rect 5742 13028 5746 13084
rect 5746 13028 5802 13084
rect 5802 13028 5806 13084
rect 5742 13024 5806 13028
rect 5822 13084 5886 13088
rect 5822 13028 5826 13084
rect 5826 13028 5882 13084
rect 5882 13028 5886 13084
rect 5822 13024 5886 13028
rect 14844 13084 14908 13088
rect 14844 13028 14848 13084
rect 14848 13028 14904 13084
rect 14904 13028 14908 13084
rect 14844 13024 14908 13028
rect 14924 13084 14988 13088
rect 14924 13028 14928 13084
rect 14928 13028 14984 13084
rect 14984 13028 14988 13084
rect 14924 13024 14988 13028
rect 15004 13084 15068 13088
rect 15004 13028 15008 13084
rect 15008 13028 15064 13084
rect 15064 13028 15068 13084
rect 15004 13024 15068 13028
rect 15084 13084 15148 13088
rect 15084 13028 15088 13084
rect 15088 13028 15144 13084
rect 15144 13028 15148 13084
rect 15084 13024 15148 13028
rect 24105 13084 24169 13088
rect 24105 13028 24109 13084
rect 24109 13028 24165 13084
rect 24165 13028 24169 13084
rect 24105 13024 24169 13028
rect 24185 13084 24249 13088
rect 24185 13028 24189 13084
rect 24189 13028 24245 13084
rect 24245 13028 24249 13084
rect 24185 13024 24249 13028
rect 24265 13084 24329 13088
rect 24265 13028 24269 13084
rect 24269 13028 24325 13084
rect 24325 13028 24329 13084
rect 24265 13024 24329 13028
rect 24345 13084 24409 13088
rect 24345 13028 24349 13084
rect 24349 13028 24405 13084
rect 24405 13028 24409 13084
rect 24345 13024 24409 13028
rect 10213 12540 10277 12544
rect 10213 12484 10217 12540
rect 10217 12484 10273 12540
rect 10273 12484 10277 12540
rect 10213 12480 10277 12484
rect 10293 12540 10357 12544
rect 10293 12484 10297 12540
rect 10297 12484 10353 12540
rect 10353 12484 10357 12540
rect 10293 12480 10357 12484
rect 10373 12540 10437 12544
rect 10373 12484 10377 12540
rect 10377 12484 10433 12540
rect 10433 12484 10437 12540
rect 10373 12480 10437 12484
rect 10453 12540 10517 12544
rect 10453 12484 10457 12540
rect 10457 12484 10513 12540
rect 10513 12484 10517 12540
rect 10453 12480 10517 12484
rect 19474 12540 19538 12544
rect 19474 12484 19478 12540
rect 19478 12484 19534 12540
rect 19534 12484 19538 12540
rect 19474 12480 19538 12484
rect 19554 12540 19618 12544
rect 19554 12484 19558 12540
rect 19558 12484 19614 12540
rect 19614 12484 19618 12540
rect 19554 12480 19618 12484
rect 19634 12540 19698 12544
rect 19634 12484 19638 12540
rect 19638 12484 19694 12540
rect 19694 12484 19698 12540
rect 19634 12480 19698 12484
rect 19714 12540 19778 12544
rect 19714 12484 19718 12540
rect 19718 12484 19774 12540
rect 19774 12484 19778 12540
rect 19714 12480 19778 12484
rect 5582 11996 5646 12000
rect 5582 11940 5586 11996
rect 5586 11940 5642 11996
rect 5642 11940 5646 11996
rect 5582 11936 5646 11940
rect 5662 11996 5726 12000
rect 5662 11940 5666 11996
rect 5666 11940 5722 11996
rect 5722 11940 5726 11996
rect 5662 11936 5726 11940
rect 5742 11996 5806 12000
rect 5742 11940 5746 11996
rect 5746 11940 5802 11996
rect 5802 11940 5806 11996
rect 5742 11936 5806 11940
rect 5822 11996 5886 12000
rect 5822 11940 5826 11996
rect 5826 11940 5882 11996
rect 5882 11940 5886 11996
rect 5822 11936 5886 11940
rect 14844 11996 14908 12000
rect 14844 11940 14848 11996
rect 14848 11940 14904 11996
rect 14904 11940 14908 11996
rect 14844 11936 14908 11940
rect 14924 11996 14988 12000
rect 14924 11940 14928 11996
rect 14928 11940 14984 11996
rect 14984 11940 14988 11996
rect 14924 11936 14988 11940
rect 15004 11996 15068 12000
rect 15004 11940 15008 11996
rect 15008 11940 15064 11996
rect 15064 11940 15068 11996
rect 15004 11936 15068 11940
rect 15084 11996 15148 12000
rect 15084 11940 15088 11996
rect 15088 11940 15144 11996
rect 15144 11940 15148 11996
rect 15084 11936 15148 11940
rect 24105 11996 24169 12000
rect 24105 11940 24109 11996
rect 24109 11940 24165 11996
rect 24165 11940 24169 11996
rect 24105 11936 24169 11940
rect 24185 11996 24249 12000
rect 24185 11940 24189 11996
rect 24189 11940 24245 11996
rect 24245 11940 24249 11996
rect 24185 11936 24249 11940
rect 24265 11996 24329 12000
rect 24265 11940 24269 11996
rect 24269 11940 24325 11996
rect 24325 11940 24329 11996
rect 24265 11936 24329 11940
rect 24345 11996 24409 12000
rect 24345 11940 24349 11996
rect 24349 11940 24405 11996
rect 24405 11940 24409 11996
rect 24345 11936 24409 11940
rect 10213 11452 10277 11456
rect 10213 11396 10217 11452
rect 10217 11396 10273 11452
rect 10273 11396 10277 11452
rect 10213 11392 10277 11396
rect 10293 11452 10357 11456
rect 10293 11396 10297 11452
rect 10297 11396 10353 11452
rect 10353 11396 10357 11452
rect 10293 11392 10357 11396
rect 10373 11452 10437 11456
rect 10373 11396 10377 11452
rect 10377 11396 10433 11452
rect 10433 11396 10437 11452
rect 10373 11392 10437 11396
rect 10453 11452 10517 11456
rect 10453 11396 10457 11452
rect 10457 11396 10513 11452
rect 10513 11396 10517 11452
rect 10453 11392 10517 11396
rect 19474 11452 19538 11456
rect 19474 11396 19478 11452
rect 19478 11396 19534 11452
rect 19534 11396 19538 11452
rect 19474 11392 19538 11396
rect 19554 11452 19618 11456
rect 19554 11396 19558 11452
rect 19558 11396 19614 11452
rect 19614 11396 19618 11452
rect 19554 11392 19618 11396
rect 19634 11452 19698 11456
rect 19634 11396 19638 11452
rect 19638 11396 19694 11452
rect 19694 11396 19698 11452
rect 19634 11392 19698 11396
rect 19714 11452 19778 11456
rect 19714 11396 19718 11452
rect 19718 11396 19774 11452
rect 19774 11396 19778 11452
rect 19714 11392 19778 11396
rect 5582 10908 5646 10912
rect 5582 10852 5586 10908
rect 5586 10852 5642 10908
rect 5642 10852 5646 10908
rect 5582 10848 5646 10852
rect 5662 10908 5726 10912
rect 5662 10852 5666 10908
rect 5666 10852 5722 10908
rect 5722 10852 5726 10908
rect 5662 10848 5726 10852
rect 5742 10908 5806 10912
rect 5742 10852 5746 10908
rect 5746 10852 5802 10908
rect 5802 10852 5806 10908
rect 5742 10848 5806 10852
rect 5822 10908 5886 10912
rect 5822 10852 5826 10908
rect 5826 10852 5882 10908
rect 5882 10852 5886 10908
rect 5822 10848 5886 10852
rect 14844 10908 14908 10912
rect 14844 10852 14848 10908
rect 14848 10852 14904 10908
rect 14904 10852 14908 10908
rect 14844 10848 14908 10852
rect 14924 10908 14988 10912
rect 14924 10852 14928 10908
rect 14928 10852 14984 10908
rect 14984 10852 14988 10908
rect 14924 10848 14988 10852
rect 15004 10908 15068 10912
rect 15004 10852 15008 10908
rect 15008 10852 15064 10908
rect 15064 10852 15068 10908
rect 15004 10848 15068 10852
rect 15084 10908 15148 10912
rect 15084 10852 15088 10908
rect 15088 10852 15144 10908
rect 15144 10852 15148 10908
rect 15084 10848 15148 10852
rect 24105 10908 24169 10912
rect 24105 10852 24109 10908
rect 24109 10852 24165 10908
rect 24165 10852 24169 10908
rect 24105 10848 24169 10852
rect 24185 10908 24249 10912
rect 24185 10852 24189 10908
rect 24189 10852 24245 10908
rect 24245 10852 24249 10908
rect 24185 10848 24249 10852
rect 24265 10908 24329 10912
rect 24265 10852 24269 10908
rect 24269 10852 24325 10908
rect 24325 10852 24329 10908
rect 24265 10848 24329 10852
rect 24345 10908 24409 10912
rect 24345 10852 24349 10908
rect 24349 10852 24405 10908
rect 24405 10852 24409 10908
rect 24345 10848 24409 10852
rect 10213 10364 10277 10368
rect 10213 10308 10217 10364
rect 10217 10308 10273 10364
rect 10273 10308 10277 10364
rect 10213 10304 10277 10308
rect 10293 10364 10357 10368
rect 10293 10308 10297 10364
rect 10297 10308 10353 10364
rect 10353 10308 10357 10364
rect 10293 10304 10357 10308
rect 10373 10364 10437 10368
rect 10373 10308 10377 10364
rect 10377 10308 10433 10364
rect 10433 10308 10437 10364
rect 10373 10304 10437 10308
rect 10453 10364 10517 10368
rect 10453 10308 10457 10364
rect 10457 10308 10513 10364
rect 10513 10308 10517 10364
rect 10453 10304 10517 10308
rect 19474 10364 19538 10368
rect 19474 10308 19478 10364
rect 19478 10308 19534 10364
rect 19534 10308 19538 10364
rect 19474 10304 19538 10308
rect 19554 10364 19618 10368
rect 19554 10308 19558 10364
rect 19558 10308 19614 10364
rect 19614 10308 19618 10364
rect 19554 10304 19618 10308
rect 19634 10364 19698 10368
rect 19634 10308 19638 10364
rect 19638 10308 19694 10364
rect 19694 10308 19698 10364
rect 19634 10304 19698 10308
rect 19714 10364 19778 10368
rect 19714 10308 19718 10364
rect 19718 10308 19774 10364
rect 19774 10308 19778 10364
rect 19714 10304 19778 10308
rect 5582 9820 5646 9824
rect 5582 9764 5586 9820
rect 5586 9764 5642 9820
rect 5642 9764 5646 9820
rect 5582 9760 5646 9764
rect 5662 9820 5726 9824
rect 5662 9764 5666 9820
rect 5666 9764 5722 9820
rect 5722 9764 5726 9820
rect 5662 9760 5726 9764
rect 5742 9820 5806 9824
rect 5742 9764 5746 9820
rect 5746 9764 5802 9820
rect 5802 9764 5806 9820
rect 5742 9760 5806 9764
rect 5822 9820 5886 9824
rect 5822 9764 5826 9820
rect 5826 9764 5882 9820
rect 5882 9764 5886 9820
rect 5822 9760 5886 9764
rect 14844 9820 14908 9824
rect 14844 9764 14848 9820
rect 14848 9764 14904 9820
rect 14904 9764 14908 9820
rect 14844 9760 14908 9764
rect 14924 9820 14988 9824
rect 14924 9764 14928 9820
rect 14928 9764 14984 9820
rect 14984 9764 14988 9820
rect 14924 9760 14988 9764
rect 15004 9820 15068 9824
rect 15004 9764 15008 9820
rect 15008 9764 15064 9820
rect 15064 9764 15068 9820
rect 15004 9760 15068 9764
rect 15084 9820 15148 9824
rect 15084 9764 15088 9820
rect 15088 9764 15144 9820
rect 15144 9764 15148 9820
rect 15084 9760 15148 9764
rect 24105 9820 24169 9824
rect 24105 9764 24109 9820
rect 24109 9764 24165 9820
rect 24165 9764 24169 9820
rect 24105 9760 24169 9764
rect 24185 9820 24249 9824
rect 24185 9764 24189 9820
rect 24189 9764 24245 9820
rect 24245 9764 24249 9820
rect 24185 9760 24249 9764
rect 24265 9820 24329 9824
rect 24265 9764 24269 9820
rect 24269 9764 24325 9820
rect 24325 9764 24329 9820
rect 24265 9760 24329 9764
rect 24345 9820 24409 9824
rect 24345 9764 24349 9820
rect 24349 9764 24405 9820
rect 24405 9764 24409 9820
rect 24345 9760 24409 9764
rect 10213 9276 10277 9280
rect 10213 9220 10217 9276
rect 10217 9220 10273 9276
rect 10273 9220 10277 9276
rect 10213 9216 10277 9220
rect 10293 9276 10357 9280
rect 10293 9220 10297 9276
rect 10297 9220 10353 9276
rect 10353 9220 10357 9276
rect 10293 9216 10357 9220
rect 10373 9276 10437 9280
rect 10373 9220 10377 9276
rect 10377 9220 10433 9276
rect 10433 9220 10437 9276
rect 10373 9216 10437 9220
rect 10453 9276 10517 9280
rect 10453 9220 10457 9276
rect 10457 9220 10513 9276
rect 10513 9220 10517 9276
rect 10453 9216 10517 9220
rect 19474 9276 19538 9280
rect 19474 9220 19478 9276
rect 19478 9220 19534 9276
rect 19534 9220 19538 9276
rect 19474 9216 19538 9220
rect 19554 9276 19618 9280
rect 19554 9220 19558 9276
rect 19558 9220 19614 9276
rect 19614 9220 19618 9276
rect 19554 9216 19618 9220
rect 19634 9276 19698 9280
rect 19634 9220 19638 9276
rect 19638 9220 19694 9276
rect 19694 9220 19698 9276
rect 19634 9216 19698 9220
rect 19714 9276 19778 9280
rect 19714 9220 19718 9276
rect 19718 9220 19774 9276
rect 19774 9220 19778 9276
rect 19714 9216 19778 9220
rect 5582 8732 5646 8736
rect 5582 8676 5586 8732
rect 5586 8676 5642 8732
rect 5642 8676 5646 8732
rect 5582 8672 5646 8676
rect 5662 8732 5726 8736
rect 5662 8676 5666 8732
rect 5666 8676 5722 8732
rect 5722 8676 5726 8732
rect 5662 8672 5726 8676
rect 5742 8732 5806 8736
rect 5742 8676 5746 8732
rect 5746 8676 5802 8732
rect 5802 8676 5806 8732
rect 5742 8672 5806 8676
rect 5822 8732 5886 8736
rect 5822 8676 5826 8732
rect 5826 8676 5882 8732
rect 5882 8676 5886 8732
rect 5822 8672 5886 8676
rect 14844 8732 14908 8736
rect 14844 8676 14848 8732
rect 14848 8676 14904 8732
rect 14904 8676 14908 8732
rect 14844 8672 14908 8676
rect 14924 8732 14988 8736
rect 14924 8676 14928 8732
rect 14928 8676 14984 8732
rect 14984 8676 14988 8732
rect 14924 8672 14988 8676
rect 15004 8732 15068 8736
rect 15004 8676 15008 8732
rect 15008 8676 15064 8732
rect 15064 8676 15068 8732
rect 15004 8672 15068 8676
rect 15084 8732 15148 8736
rect 15084 8676 15088 8732
rect 15088 8676 15144 8732
rect 15144 8676 15148 8732
rect 15084 8672 15148 8676
rect 24105 8732 24169 8736
rect 24105 8676 24109 8732
rect 24109 8676 24165 8732
rect 24165 8676 24169 8732
rect 24105 8672 24169 8676
rect 24185 8732 24249 8736
rect 24185 8676 24189 8732
rect 24189 8676 24245 8732
rect 24245 8676 24249 8732
rect 24185 8672 24249 8676
rect 24265 8732 24329 8736
rect 24265 8676 24269 8732
rect 24269 8676 24325 8732
rect 24325 8676 24329 8732
rect 24265 8672 24329 8676
rect 24345 8732 24409 8736
rect 24345 8676 24349 8732
rect 24349 8676 24405 8732
rect 24405 8676 24409 8732
rect 24345 8672 24409 8676
rect 10213 8188 10277 8192
rect 10213 8132 10217 8188
rect 10217 8132 10273 8188
rect 10273 8132 10277 8188
rect 10213 8128 10277 8132
rect 10293 8188 10357 8192
rect 10293 8132 10297 8188
rect 10297 8132 10353 8188
rect 10353 8132 10357 8188
rect 10293 8128 10357 8132
rect 10373 8188 10437 8192
rect 10373 8132 10377 8188
rect 10377 8132 10433 8188
rect 10433 8132 10437 8188
rect 10373 8128 10437 8132
rect 10453 8188 10517 8192
rect 10453 8132 10457 8188
rect 10457 8132 10513 8188
rect 10513 8132 10517 8188
rect 10453 8128 10517 8132
rect 19474 8188 19538 8192
rect 19474 8132 19478 8188
rect 19478 8132 19534 8188
rect 19534 8132 19538 8188
rect 19474 8128 19538 8132
rect 19554 8188 19618 8192
rect 19554 8132 19558 8188
rect 19558 8132 19614 8188
rect 19614 8132 19618 8188
rect 19554 8128 19618 8132
rect 19634 8188 19698 8192
rect 19634 8132 19638 8188
rect 19638 8132 19694 8188
rect 19694 8132 19698 8188
rect 19634 8128 19698 8132
rect 19714 8188 19778 8192
rect 19714 8132 19718 8188
rect 19718 8132 19774 8188
rect 19774 8132 19778 8188
rect 19714 8128 19778 8132
rect 5582 7644 5646 7648
rect 5582 7588 5586 7644
rect 5586 7588 5642 7644
rect 5642 7588 5646 7644
rect 5582 7584 5646 7588
rect 5662 7644 5726 7648
rect 5662 7588 5666 7644
rect 5666 7588 5722 7644
rect 5722 7588 5726 7644
rect 5662 7584 5726 7588
rect 5742 7644 5806 7648
rect 5742 7588 5746 7644
rect 5746 7588 5802 7644
rect 5802 7588 5806 7644
rect 5742 7584 5806 7588
rect 5822 7644 5886 7648
rect 5822 7588 5826 7644
rect 5826 7588 5882 7644
rect 5882 7588 5886 7644
rect 5822 7584 5886 7588
rect 14844 7644 14908 7648
rect 14844 7588 14848 7644
rect 14848 7588 14904 7644
rect 14904 7588 14908 7644
rect 14844 7584 14908 7588
rect 14924 7644 14988 7648
rect 14924 7588 14928 7644
rect 14928 7588 14984 7644
rect 14984 7588 14988 7644
rect 14924 7584 14988 7588
rect 15004 7644 15068 7648
rect 15004 7588 15008 7644
rect 15008 7588 15064 7644
rect 15064 7588 15068 7644
rect 15004 7584 15068 7588
rect 15084 7644 15148 7648
rect 15084 7588 15088 7644
rect 15088 7588 15144 7644
rect 15144 7588 15148 7644
rect 15084 7584 15148 7588
rect 24105 7644 24169 7648
rect 24105 7588 24109 7644
rect 24109 7588 24165 7644
rect 24165 7588 24169 7644
rect 24105 7584 24169 7588
rect 24185 7644 24249 7648
rect 24185 7588 24189 7644
rect 24189 7588 24245 7644
rect 24245 7588 24249 7644
rect 24185 7584 24249 7588
rect 24265 7644 24329 7648
rect 24265 7588 24269 7644
rect 24269 7588 24325 7644
rect 24325 7588 24329 7644
rect 24265 7584 24329 7588
rect 24345 7644 24409 7648
rect 24345 7588 24349 7644
rect 24349 7588 24405 7644
rect 24405 7588 24409 7644
rect 24345 7584 24409 7588
rect 10213 7100 10277 7104
rect 10213 7044 10217 7100
rect 10217 7044 10273 7100
rect 10273 7044 10277 7100
rect 10213 7040 10277 7044
rect 10293 7100 10357 7104
rect 10293 7044 10297 7100
rect 10297 7044 10353 7100
rect 10353 7044 10357 7100
rect 10293 7040 10357 7044
rect 10373 7100 10437 7104
rect 10373 7044 10377 7100
rect 10377 7044 10433 7100
rect 10433 7044 10437 7100
rect 10373 7040 10437 7044
rect 10453 7100 10517 7104
rect 10453 7044 10457 7100
rect 10457 7044 10513 7100
rect 10513 7044 10517 7100
rect 10453 7040 10517 7044
rect 19474 7100 19538 7104
rect 19474 7044 19478 7100
rect 19478 7044 19534 7100
rect 19534 7044 19538 7100
rect 19474 7040 19538 7044
rect 19554 7100 19618 7104
rect 19554 7044 19558 7100
rect 19558 7044 19614 7100
rect 19614 7044 19618 7100
rect 19554 7040 19618 7044
rect 19634 7100 19698 7104
rect 19634 7044 19638 7100
rect 19638 7044 19694 7100
rect 19694 7044 19698 7100
rect 19634 7040 19698 7044
rect 19714 7100 19778 7104
rect 19714 7044 19718 7100
rect 19718 7044 19774 7100
rect 19774 7044 19778 7100
rect 19714 7040 19778 7044
rect 5582 6556 5646 6560
rect 5582 6500 5586 6556
rect 5586 6500 5642 6556
rect 5642 6500 5646 6556
rect 5582 6496 5646 6500
rect 5662 6556 5726 6560
rect 5662 6500 5666 6556
rect 5666 6500 5722 6556
rect 5722 6500 5726 6556
rect 5662 6496 5726 6500
rect 5742 6556 5806 6560
rect 5742 6500 5746 6556
rect 5746 6500 5802 6556
rect 5802 6500 5806 6556
rect 5742 6496 5806 6500
rect 5822 6556 5886 6560
rect 5822 6500 5826 6556
rect 5826 6500 5882 6556
rect 5882 6500 5886 6556
rect 5822 6496 5886 6500
rect 14844 6556 14908 6560
rect 14844 6500 14848 6556
rect 14848 6500 14904 6556
rect 14904 6500 14908 6556
rect 14844 6496 14908 6500
rect 14924 6556 14988 6560
rect 14924 6500 14928 6556
rect 14928 6500 14984 6556
rect 14984 6500 14988 6556
rect 14924 6496 14988 6500
rect 15004 6556 15068 6560
rect 15004 6500 15008 6556
rect 15008 6500 15064 6556
rect 15064 6500 15068 6556
rect 15004 6496 15068 6500
rect 15084 6556 15148 6560
rect 15084 6500 15088 6556
rect 15088 6500 15144 6556
rect 15144 6500 15148 6556
rect 15084 6496 15148 6500
rect 24105 6556 24169 6560
rect 24105 6500 24109 6556
rect 24109 6500 24165 6556
rect 24165 6500 24169 6556
rect 24105 6496 24169 6500
rect 24185 6556 24249 6560
rect 24185 6500 24189 6556
rect 24189 6500 24245 6556
rect 24245 6500 24249 6556
rect 24185 6496 24249 6500
rect 24265 6556 24329 6560
rect 24265 6500 24269 6556
rect 24269 6500 24325 6556
rect 24325 6500 24329 6556
rect 24265 6496 24329 6500
rect 24345 6556 24409 6560
rect 24345 6500 24349 6556
rect 24349 6500 24405 6556
rect 24405 6500 24409 6556
rect 24345 6496 24409 6500
rect 10213 6012 10277 6016
rect 10213 5956 10217 6012
rect 10217 5956 10273 6012
rect 10273 5956 10277 6012
rect 10213 5952 10277 5956
rect 10293 6012 10357 6016
rect 10293 5956 10297 6012
rect 10297 5956 10353 6012
rect 10353 5956 10357 6012
rect 10293 5952 10357 5956
rect 10373 6012 10437 6016
rect 10373 5956 10377 6012
rect 10377 5956 10433 6012
rect 10433 5956 10437 6012
rect 10373 5952 10437 5956
rect 10453 6012 10517 6016
rect 10453 5956 10457 6012
rect 10457 5956 10513 6012
rect 10513 5956 10517 6012
rect 10453 5952 10517 5956
rect 19474 6012 19538 6016
rect 19474 5956 19478 6012
rect 19478 5956 19534 6012
rect 19534 5956 19538 6012
rect 19474 5952 19538 5956
rect 19554 6012 19618 6016
rect 19554 5956 19558 6012
rect 19558 5956 19614 6012
rect 19614 5956 19618 6012
rect 19554 5952 19618 5956
rect 19634 6012 19698 6016
rect 19634 5956 19638 6012
rect 19638 5956 19694 6012
rect 19694 5956 19698 6012
rect 19634 5952 19698 5956
rect 19714 6012 19778 6016
rect 19714 5956 19718 6012
rect 19718 5956 19774 6012
rect 19774 5956 19778 6012
rect 19714 5952 19778 5956
rect 5582 5468 5646 5472
rect 5582 5412 5586 5468
rect 5586 5412 5642 5468
rect 5642 5412 5646 5468
rect 5582 5408 5646 5412
rect 5662 5468 5726 5472
rect 5662 5412 5666 5468
rect 5666 5412 5722 5468
rect 5722 5412 5726 5468
rect 5662 5408 5726 5412
rect 5742 5468 5806 5472
rect 5742 5412 5746 5468
rect 5746 5412 5802 5468
rect 5802 5412 5806 5468
rect 5742 5408 5806 5412
rect 5822 5468 5886 5472
rect 5822 5412 5826 5468
rect 5826 5412 5882 5468
rect 5882 5412 5886 5468
rect 5822 5408 5886 5412
rect 14844 5468 14908 5472
rect 14844 5412 14848 5468
rect 14848 5412 14904 5468
rect 14904 5412 14908 5468
rect 14844 5408 14908 5412
rect 14924 5468 14988 5472
rect 14924 5412 14928 5468
rect 14928 5412 14984 5468
rect 14984 5412 14988 5468
rect 14924 5408 14988 5412
rect 15004 5468 15068 5472
rect 15004 5412 15008 5468
rect 15008 5412 15064 5468
rect 15064 5412 15068 5468
rect 15004 5408 15068 5412
rect 15084 5468 15148 5472
rect 15084 5412 15088 5468
rect 15088 5412 15144 5468
rect 15144 5412 15148 5468
rect 15084 5408 15148 5412
rect 24105 5468 24169 5472
rect 24105 5412 24109 5468
rect 24109 5412 24165 5468
rect 24165 5412 24169 5468
rect 24105 5408 24169 5412
rect 24185 5468 24249 5472
rect 24185 5412 24189 5468
rect 24189 5412 24245 5468
rect 24245 5412 24249 5468
rect 24185 5408 24249 5412
rect 24265 5468 24329 5472
rect 24265 5412 24269 5468
rect 24269 5412 24325 5468
rect 24325 5412 24329 5468
rect 24265 5408 24329 5412
rect 24345 5468 24409 5472
rect 24345 5412 24349 5468
rect 24349 5412 24405 5468
rect 24405 5412 24409 5468
rect 24345 5408 24409 5412
rect 10213 4924 10277 4928
rect 10213 4868 10217 4924
rect 10217 4868 10273 4924
rect 10273 4868 10277 4924
rect 10213 4864 10277 4868
rect 10293 4924 10357 4928
rect 10293 4868 10297 4924
rect 10297 4868 10353 4924
rect 10353 4868 10357 4924
rect 10293 4864 10357 4868
rect 10373 4924 10437 4928
rect 10373 4868 10377 4924
rect 10377 4868 10433 4924
rect 10433 4868 10437 4924
rect 10373 4864 10437 4868
rect 10453 4924 10517 4928
rect 10453 4868 10457 4924
rect 10457 4868 10513 4924
rect 10513 4868 10517 4924
rect 10453 4864 10517 4868
rect 19474 4924 19538 4928
rect 19474 4868 19478 4924
rect 19478 4868 19534 4924
rect 19534 4868 19538 4924
rect 19474 4864 19538 4868
rect 19554 4924 19618 4928
rect 19554 4868 19558 4924
rect 19558 4868 19614 4924
rect 19614 4868 19618 4924
rect 19554 4864 19618 4868
rect 19634 4924 19698 4928
rect 19634 4868 19638 4924
rect 19638 4868 19694 4924
rect 19694 4868 19698 4924
rect 19634 4864 19698 4868
rect 19714 4924 19778 4928
rect 19714 4868 19718 4924
rect 19718 4868 19774 4924
rect 19774 4868 19778 4924
rect 19714 4864 19778 4868
rect 5582 4380 5646 4384
rect 5582 4324 5586 4380
rect 5586 4324 5642 4380
rect 5642 4324 5646 4380
rect 5582 4320 5646 4324
rect 5662 4380 5726 4384
rect 5662 4324 5666 4380
rect 5666 4324 5722 4380
rect 5722 4324 5726 4380
rect 5662 4320 5726 4324
rect 5742 4380 5806 4384
rect 5742 4324 5746 4380
rect 5746 4324 5802 4380
rect 5802 4324 5806 4380
rect 5742 4320 5806 4324
rect 5822 4380 5886 4384
rect 5822 4324 5826 4380
rect 5826 4324 5882 4380
rect 5882 4324 5886 4380
rect 5822 4320 5886 4324
rect 14844 4380 14908 4384
rect 14844 4324 14848 4380
rect 14848 4324 14904 4380
rect 14904 4324 14908 4380
rect 14844 4320 14908 4324
rect 14924 4380 14988 4384
rect 14924 4324 14928 4380
rect 14928 4324 14984 4380
rect 14984 4324 14988 4380
rect 14924 4320 14988 4324
rect 15004 4380 15068 4384
rect 15004 4324 15008 4380
rect 15008 4324 15064 4380
rect 15064 4324 15068 4380
rect 15004 4320 15068 4324
rect 15084 4380 15148 4384
rect 15084 4324 15088 4380
rect 15088 4324 15144 4380
rect 15144 4324 15148 4380
rect 15084 4320 15148 4324
rect 24105 4380 24169 4384
rect 24105 4324 24109 4380
rect 24109 4324 24165 4380
rect 24165 4324 24169 4380
rect 24105 4320 24169 4324
rect 24185 4380 24249 4384
rect 24185 4324 24189 4380
rect 24189 4324 24245 4380
rect 24245 4324 24249 4380
rect 24185 4320 24249 4324
rect 24265 4380 24329 4384
rect 24265 4324 24269 4380
rect 24269 4324 24325 4380
rect 24325 4324 24329 4380
rect 24265 4320 24329 4324
rect 24345 4380 24409 4384
rect 24345 4324 24349 4380
rect 24349 4324 24405 4380
rect 24405 4324 24409 4380
rect 24345 4320 24409 4324
rect 10213 3836 10277 3840
rect 10213 3780 10217 3836
rect 10217 3780 10273 3836
rect 10273 3780 10277 3836
rect 10213 3776 10277 3780
rect 10293 3836 10357 3840
rect 10293 3780 10297 3836
rect 10297 3780 10353 3836
rect 10353 3780 10357 3836
rect 10293 3776 10357 3780
rect 10373 3836 10437 3840
rect 10373 3780 10377 3836
rect 10377 3780 10433 3836
rect 10433 3780 10437 3836
rect 10373 3776 10437 3780
rect 10453 3836 10517 3840
rect 10453 3780 10457 3836
rect 10457 3780 10513 3836
rect 10513 3780 10517 3836
rect 10453 3776 10517 3780
rect 19474 3836 19538 3840
rect 19474 3780 19478 3836
rect 19478 3780 19534 3836
rect 19534 3780 19538 3836
rect 19474 3776 19538 3780
rect 19554 3836 19618 3840
rect 19554 3780 19558 3836
rect 19558 3780 19614 3836
rect 19614 3780 19618 3836
rect 19554 3776 19618 3780
rect 19634 3836 19698 3840
rect 19634 3780 19638 3836
rect 19638 3780 19694 3836
rect 19694 3780 19698 3836
rect 19634 3776 19698 3780
rect 19714 3836 19778 3840
rect 19714 3780 19718 3836
rect 19718 3780 19774 3836
rect 19774 3780 19778 3836
rect 19714 3776 19778 3780
rect 5582 3292 5646 3296
rect 5582 3236 5586 3292
rect 5586 3236 5642 3292
rect 5642 3236 5646 3292
rect 5582 3232 5646 3236
rect 5662 3292 5726 3296
rect 5662 3236 5666 3292
rect 5666 3236 5722 3292
rect 5722 3236 5726 3292
rect 5662 3232 5726 3236
rect 5742 3292 5806 3296
rect 5742 3236 5746 3292
rect 5746 3236 5802 3292
rect 5802 3236 5806 3292
rect 5742 3232 5806 3236
rect 5822 3292 5886 3296
rect 5822 3236 5826 3292
rect 5826 3236 5882 3292
rect 5882 3236 5886 3292
rect 5822 3232 5886 3236
rect 14844 3292 14908 3296
rect 14844 3236 14848 3292
rect 14848 3236 14904 3292
rect 14904 3236 14908 3292
rect 14844 3232 14908 3236
rect 14924 3292 14988 3296
rect 14924 3236 14928 3292
rect 14928 3236 14984 3292
rect 14984 3236 14988 3292
rect 14924 3232 14988 3236
rect 15004 3292 15068 3296
rect 15004 3236 15008 3292
rect 15008 3236 15064 3292
rect 15064 3236 15068 3292
rect 15004 3232 15068 3236
rect 15084 3292 15148 3296
rect 15084 3236 15088 3292
rect 15088 3236 15144 3292
rect 15144 3236 15148 3292
rect 15084 3232 15148 3236
rect 24105 3292 24169 3296
rect 24105 3236 24109 3292
rect 24109 3236 24165 3292
rect 24165 3236 24169 3292
rect 24105 3232 24169 3236
rect 24185 3292 24249 3296
rect 24185 3236 24189 3292
rect 24189 3236 24245 3292
rect 24245 3236 24249 3292
rect 24185 3232 24249 3236
rect 24265 3292 24329 3296
rect 24265 3236 24269 3292
rect 24269 3236 24325 3292
rect 24325 3236 24329 3292
rect 24265 3232 24329 3236
rect 24345 3292 24409 3296
rect 24345 3236 24349 3292
rect 24349 3236 24405 3292
rect 24405 3236 24409 3292
rect 24345 3232 24409 3236
rect 10213 2748 10277 2752
rect 10213 2692 10217 2748
rect 10217 2692 10273 2748
rect 10273 2692 10277 2748
rect 10213 2688 10277 2692
rect 10293 2748 10357 2752
rect 10293 2692 10297 2748
rect 10297 2692 10353 2748
rect 10353 2692 10357 2748
rect 10293 2688 10357 2692
rect 10373 2748 10437 2752
rect 10373 2692 10377 2748
rect 10377 2692 10433 2748
rect 10433 2692 10437 2748
rect 10373 2688 10437 2692
rect 10453 2748 10517 2752
rect 10453 2692 10457 2748
rect 10457 2692 10513 2748
rect 10513 2692 10517 2748
rect 10453 2688 10517 2692
rect 19474 2748 19538 2752
rect 19474 2692 19478 2748
rect 19478 2692 19534 2748
rect 19534 2692 19538 2748
rect 19474 2688 19538 2692
rect 19554 2748 19618 2752
rect 19554 2692 19558 2748
rect 19558 2692 19614 2748
rect 19614 2692 19618 2748
rect 19554 2688 19618 2692
rect 19634 2748 19698 2752
rect 19634 2692 19638 2748
rect 19638 2692 19694 2748
rect 19694 2692 19698 2748
rect 19634 2688 19698 2692
rect 19714 2748 19778 2752
rect 19714 2692 19718 2748
rect 19718 2692 19774 2748
rect 19774 2692 19778 2748
rect 19714 2688 19778 2692
rect 5582 2204 5646 2208
rect 5582 2148 5586 2204
rect 5586 2148 5642 2204
rect 5642 2148 5646 2204
rect 5582 2144 5646 2148
rect 5662 2204 5726 2208
rect 5662 2148 5666 2204
rect 5666 2148 5722 2204
rect 5722 2148 5726 2204
rect 5662 2144 5726 2148
rect 5742 2204 5806 2208
rect 5742 2148 5746 2204
rect 5746 2148 5802 2204
rect 5802 2148 5806 2204
rect 5742 2144 5806 2148
rect 5822 2204 5886 2208
rect 5822 2148 5826 2204
rect 5826 2148 5882 2204
rect 5882 2148 5886 2204
rect 5822 2144 5886 2148
rect 14844 2204 14908 2208
rect 14844 2148 14848 2204
rect 14848 2148 14904 2204
rect 14904 2148 14908 2204
rect 14844 2144 14908 2148
rect 14924 2204 14988 2208
rect 14924 2148 14928 2204
rect 14928 2148 14984 2204
rect 14984 2148 14988 2204
rect 14924 2144 14988 2148
rect 15004 2204 15068 2208
rect 15004 2148 15008 2204
rect 15008 2148 15064 2204
rect 15064 2148 15068 2204
rect 15004 2144 15068 2148
rect 15084 2204 15148 2208
rect 15084 2148 15088 2204
rect 15088 2148 15144 2204
rect 15144 2148 15148 2204
rect 15084 2144 15148 2148
rect 24105 2204 24169 2208
rect 24105 2148 24109 2204
rect 24109 2148 24165 2204
rect 24165 2148 24169 2204
rect 24105 2144 24169 2148
rect 24185 2204 24249 2208
rect 24185 2148 24189 2204
rect 24189 2148 24245 2204
rect 24245 2148 24249 2204
rect 24185 2144 24249 2148
rect 24265 2204 24329 2208
rect 24265 2148 24269 2204
rect 24269 2148 24325 2204
rect 24325 2148 24329 2204
rect 24265 2144 24329 2148
rect 24345 2204 24409 2208
rect 24345 2148 24349 2204
rect 24349 2148 24405 2204
rect 24405 2148 24409 2204
rect 24345 2144 24409 2148
<< metal4 >>
rect 5574 29408 5895 29968
rect 5574 29344 5582 29408
rect 5646 29344 5662 29408
rect 5726 29344 5742 29408
rect 5806 29344 5822 29408
rect 5886 29344 5895 29408
rect 5574 28320 5895 29344
rect 5574 28256 5582 28320
rect 5646 28256 5662 28320
rect 5726 28256 5742 28320
rect 5806 28256 5822 28320
rect 5886 28256 5895 28320
rect 5574 27232 5895 28256
rect 5574 27168 5582 27232
rect 5646 27168 5662 27232
rect 5726 27168 5742 27232
rect 5806 27168 5822 27232
rect 5886 27168 5895 27232
rect 5574 26144 5895 27168
rect 5574 26080 5582 26144
rect 5646 26080 5662 26144
rect 5726 26080 5742 26144
rect 5806 26080 5822 26144
rect 5886 26080 5895 26144
rect 5574 25366 5895 26080
rect 5574 25130 5616 25366
rect 5852 25130 5895 25366
rect 5574 25056 5895 25130
rect 5574 24992 5582 25056
rect 5646 24992 5662 25056
rect 5726 24992 5742 25056
rect 5806 24992 5822 25056
rect 5886 24992 5895 25056
rect 5574 23968 5895 24992
rect 5574 23904 5582 23968
rect 5646 23904 5662 23968
rect 5726 23904 5742 23968
rect 5806 23904 5822 23968
rect 5886 23904 5895 23968
rect 5574 22880 5895 23904
rect 5574 22816 5582 22880
rect 5646 22816 5662 22880
rect 5726 22816 5742 22880
rect 5806 22816 5822 22880
rect 5886 22816 5895 22880
rect 5574 21792 5895 22816
rect 5574 21728 5582 21792
rect 5646 21728 5662 21792
rect 5726 21728 5742 21792
rect 5806 21728 5822 21792
rect 5886 21728 5895 21792
rect 5574 20704 5895 21728
rect 5574 20640 5582 20704
rect 5646 20640 5662 20704
rect 5726 20640 5742 20704
rect 5806 20640 5822 20704
rect 5886 20640 5895 20704
rect 5574 19616 5895 20640
rect 5574 19552 5582 19616
rect 5646 19552 5662 19616
rect 5726 19552 5742 19616
rect 5806 19552 5822 19616
rect 5886 19552 5895 19616
rect 5574 18528 5895 19552
rect 5574 18464 5582 18528
rect 5646 18464 5662 18528
rect 5726 18464 5742 18528
rect 5806 18464 5822 18528
rect 5886 18464 5895 18528
rect 5574 17440 5895 18464
rect 5574 17376 5582 17440
rect 5646 17376 5662 17440
rect 5726 17376 5742 17440
rect 5806 17376 5822 17440
rect 5886 17376 5895 17440
rect 5574 16352 5895 17376
rect 5574 16288 5582 16352
rect 5646 16288 5662 16352
rect 5726 16288 5742 16352
rect 5806 16288 5822 16352
rect 5886 16288 5895 16352
rect 5574 16118 5895 16288
rect 5574 15882 5616 16118
rect 5852 15882 5895 16118
rect 5574 15264 5895 15882
rect 5574 15200 5582 15264
rect 5646 15200 5662 15264
rect 5726 15200 5742 15264
rect 5806 15200 5822 15264
rect 5886 15200 5895 15264
rect 5574 14176 5895 15200
rect 5574 14112 5582 14176
rect 5646 14112 5662 14176
rect 5726 14112 5742 14176
rect 5806 14112 5822 14176
rect 5886 14112 5895 14176
rect 5574 13088 5895 14112
rect 5574 13024 5582 13088
rect 5646 13024 5662 13088
rect 5726 13024 5742 13088
rect 5806 13024 5822 13088
rect 5886 13024 5895 13088
rect 5574 12000 5895 13024
rect 5574 11936 5582 12000
rect 5646 11936 5662 12000
rect 5726 11936 5742 12000
rect 5806 11936 5822 12000
rect 5886 11936 5895 12000
rect 5574 10912 5895 11936
rect 5574 10848 5582 10912
rect 5646 10848 5662 10912
rect 5726 10848 5742 10912
rect 5806 10848 5822 10912
rect 5886 10848 5895 10912
rect 5574 9824 5895 10848
rect 5574 9760 5582 9824
rect 5646 9760 5662 9824
rect 5726 9760 5742 9824
rect 5806 9760 5822 9824
rect 5886 9760 5895 9824
rect 5574 8736 5895 9760
rect 5574 8672 5582 8736
rect 5646 8672 5662 8736
rect 5726 8672 5742 8736
rect 5806 8672 5822 8736
rect 5886 8672 5895 8736
rect 5574 7648 5895 8672
rect 5574 7584 5582 7648
rect 5646 7584 5662 7648
rect 5726 7584 5742 7648
rect 5806 7584 5822 7648
rect 5886 7584 5895 7648
rect 5574 6870 5895 7584
rect 5574 6634 5616 6870
rect 5852 6634 5895 6870
rect 5574 6560 5895 6634
rect 5574 6496 5582 6560
rect 5646 6496 5662 6560
rect 5726 6496 5742 6560
rect 5806 6496 5822 6560
rect 5886 6496 5895 6560
rect 5574 5472 5895 6496
rect 5574 5408 5582 5472
rect 5646 5408 5662 5472
rect 5726 5408 5742 5472
rect 5806 5408 5822 5472
rect 5886 5408 5895 5472
rect 5574 4384 5895 5408
rect 5574 4320 5582 4384
rect 5646 4320 5662 4384
rect 5726 4320 5742 4384
rect 5806 4320 5822 4384
rect 5886 4320 5895 4384
rect 5574 3296 5895 4320
rect 5574 3232 5582 3296
rect 5646 3232 5662 3296
rect 5726 3232 5742 3296
rect 5806 3232 5822 3296
rect 5886 3232 5895 3296
rect 5574 2208 5895 3232
rect 5574 2144 5582 2208
rect 5646 2144 5662 2208
rect 5726 2144 5742 2208
rect 5806 2144 5822 2208
rect 5886 2144 5895 2208
rect 5574 2128 5895 2144
rect 10205 29952 10525 29968
rect 10205 29888 10213 29952
rect 10277 29888 10293 29952
rect 10357 29888 10373 29952
rect 10437 29888 10453 29952
rect 10517 29888 10525 29952
rect 10205 28864 10525 29888
rect 10205 28800 10213 28864
rect 10277 28800 10293 28864
rect 10357 28800 10373 28864
rect 10437 28800 10453 28864
rect 10517 28800 10525 28864
rect 10205 27776 10525 28800
rect 10205 27712 10213 27776
rect 10277 27712 10293 27776
rect 10357 27712 10373 27776
rect 10437 27712 10453 27776
rect 10517 27712 10525 27776
rect 10205 26688 10525 27712
rect 10205 26624 10213 26688
rect 10277 26624 10293 26688
rect 10357 26624 10373 26688
rect 10437 26624 10453 26688
rect 10517 26624 10525 26688
rect 10205 25600 10525 26624
rect 10205 25536 10213 25600
rect 10277 25536 10293 25600
rect 10357 25536 10373 25600
rect 10437 25536 10453 25600
rect 10517 25536 10525 25600
rect 10205 24512 10525 25536
rect 10205 24448 10213 24512
rect 10277 24448 10293 24512
rect 10357 24448 10373 24512
rect 10437 24448 10453 24512
rect 10517 24448 10525 24512
rect 10205 23424 10525 24448
rect 10205 23360 10213 23424
rect 10277 23360 10293 23424
rect 10357 23360 10373 23424
rect 10437 23360 10453 23424
rect 10517 23360 10525 23424
rect 10205 22336 10525 23360
rect 10205 22272 10213 22336
rect 10277 22272 10293 22336
rect 10357 22272 10373 22336
rect 10437 22272 10453 22336
rect 10517 22272 10525 22336
rect 10205 21248 10525 22272
rect 10205 21184 10213 21248
rect 10277 21184 10293 21248
rect 10357 21184 10373 21248
rect 10437 21184 10453 21248
rect 10517 21184 10525 21248
rect 10205 20742 10525 21184
rect 10205 20506 10247 20742
rect 10483 20506 10525 20742
rect 10205 20160 10525 20506
rect 10205 20096 10213 20160
rect 10277 20096 10293 20160
rect 10357 20096 10373 20160
rect 10437 20096 10453 20160
rect 10517 20096 10525 20160
rect 10205 19072 10525 20096
rect 10205 19008 10213 19072
rect 10277 19008 10293 19072
rect 10357 19008 10373 19072
rect 10437 19008 10453 19072
rect 10517 19008 10525 19072
rect 10205 17984 10525 19008
rect 10205 17920 10213 17984
rect 10277 17920 10293 17984
rect 10357 17920 10373 17984
rect 10437 17920 10453 17984
rect 10517 17920 10525 17984
rect 10205 16896 10525 17920
rect 10205 16832 10213 16896
rect 10277 16832 10293 16896
rect 10357 16832 10373 16896
rect 10437 16832 10453 16896
rect 10517 16832 10525 16896
rect 10205 15808 10525 16832
rect 10205 15744 10213 15808
rect 10277 15744 10293 15808
rect 10357 15744 10373 15808
rect 10437 15744 10453 15808
rect 10517 15744 10525 15808
rect 10205 14720 10525 15744
rect 10205 14656 10213 14720
rect 10277 14656 10293 14720
rect 10357 14656 10373 14720
rect 10437 14656 10453 14720
rect 10517 14656 10525 14720
rect 10205 13632 10525 14656
rect 10205 13568 10213 13632
rect 10277 13568 10293 13632
rect 10357 13568 10373 13632
rect 10437 13568 10453 13632
rect 10517 13568 10525 13632
rect 10205 12544 10525 13568
rect 10205 12480 10213 12544
rect 10277 12480 10293 12544
rect 10357 12480 10373 12544
rect 10437 12480 10453 12544
rect 10517 12480 10525 12544
rect 10205 11494 10525 12480
rect 10205 11456 10247 11494
rect 10483 11456 10525 11494
rect 10205 11392 10213 11456
rect 10517 11392 10525 11456
rect 10205 11258 10247 11392
rect 10483 11258 10525 11392
rect 10205 10368 10525 11258
rect 10205 10304 10213 10368
rect 10277 10304 10293 10368
rect 10357 10304 10373 10368
rect 10437 10304 10453 10368
rect 10517 10304 10525 10368
rect 10205 9280 10525 10304
rect 10205 9216 10213 9280
rect 10277 9216 10293 9280
rect 10357 9216 10373 9280
rect 10437 9216 10453 9280
rect 10517 9216 10525 9280
rect 10205 8192 10525 9216
rect 10205 8128 10213 8192
rect 10277 8128 10293 8192
rect 10357 8128 10373 8192
rect 10437 8128 10453 8192
rect 10517 8128 10525 8192
rect 10205 7104 10525 8128
rect 10205 7040 10213 7104
rect 10277 7040 10293 7104
rect 10357 7040 10373 7104
rect 10437 7040 10453 7104
rect 10517 7040 10525 7104
rect 10205 6016 10525 7040
rect 10205 5952 10213 6016
rect 10277 5952 10293 6016
rect 10357 5952 10373 6016
rect 10437 5952 10453 6016
rect 10517 5952 10525 6016
rect 10205 4928 10525 5952
rect 10205 4864 10213 4928
rect 10277 4864 10293 4928
rect 10357 4864 10373 4928
rect 10437 4864 10453 4928
rect 10517 4864 10525 4928
rect 10205 3840 10525 4864
rect 10205 3776 10213 3840
rect 10277 3776 10293 3840
rect 10357 3776 10373 3840
rect 10437 3776 10453 3840
rect 10517 3776 10525 3840
rect 10205 2752 10525 3776
rect 10205 2688 10213 2752
rect 10277 2688 10293 2752
rect 10357 2688 10373 2752
rect 10437 2688 10453 2752
rect 10517 2688 10525 2752
rect 10205 2128 10525 2688
rect 14836 29408 15156 29968
rect 14836 29344 14844 29408
rect 14908 29344 14924 29408
rect 14988 29344 15004 29408
rect 15068 29344 15084 29408
rect 15148 29344 15156 29408
rect 14836 28320 15156 29344
rect 14836 28256 14844 28320
rect 14908 28256 14924 28320
rect 14988 28256 15004 28320
rect 15068 28256 15084 28320
rect 15148 28256 15156 28320
rect 14836 27232 15156 28256
rect 14836 27168 14844 27232
rect 14908 27168 14924 27232
rect 14988 27168 15004 27232
rect 15068 27168 15084 27232
rect 15148 27168 15156 27232
rect 14836 26144 15156 27168
rect 14836 26080 14844 26144
rect 14908 26080 14924 26144
rect 14988 26080 15004 26144
rect 15068 26080 15084 26144
rect 15148 26080 15156 26144
rect 14836 25366 15156 26080
rect 14836 25130 14878 25366
rect 15114 25130 15156 25366
rect 14836 25056 15156 25130
rect 14836 24992 14844 25056
rect 14908 24992 14924 25056
rect 14988 24992 15004 25056
rect 15068 24992 15084 25056
rect 15148 24992 15156 25056
rect 14836 23968 15156 24992
rect 14836 23904 14844 23968
rect 14908 23904 14924 23968
rect 14988 23904 15004 23968
rect 15068 23904 15084 23968
rect 15148 23904 15156 23968
rect 14836 22880 15156 23904
rect 14836 22816 14844 22880
rect 14908 22816 14924 22880
rect 14988 22816 15004 22880
rect 15068 22816 15084 22880
rect 15148 22816 15156 22880
rect 14836 21792 15156 22816
rect 14836 21728 14844 21792
rect 14908 21728 14924 21792
rect 14988 21728 15004 21792
rect 15068 21728 15084 21792
rect 15148 21728 15156 21792
rect 14836 20704 15156 21728
rect 14836 20640 14844 20704
rect 14908 20640 14924 20704
rect 14988 20640 15004 20704
rect 15068 20640 15084 20704
rect 15148 20640 15156 20704
rect 14836 19616 15156 20640
rect 14836 19552 14844 19616
rect 14908 19552 14924 19616
rect 14988 19552 15004 19616
rect 15068 19552 15084 19616
rect 15148 19552 15156 19616
rect 14836 18528 15156 19552
rect 14836 18464 14844 18528
rect 14908 18464 14924 18528
rect 14988 18464 15004 18528
rect 15068 18464 15084 18528
rect 15148 18464 15156 18528
rect 14836 17440 15156 18464
rect 14836 17376 14844 17440
rect 14908 17376 14924 17440
rect 14988 17376 15004 17440
rect 15068 17376 15084 17440
rect 15148 17376 15156 17440
rect 14836 16352 15156 17376
rect 14836 16288 14844 16352
rect 14908 16288 14924 16352
rect 14988 16288 15004 16352
rect 15068 16288 15084 16352
rect 15148 16288 15156 16352
rect 14836 16118 15156 16288
rect 14836 15882 14878 16118
rect 15114 15882 15156 16118
rect 14836 15264 15156 15882
rect 14836 15200 14844 15264
rect 14908 15200 14924 15264
rect 14988 15200 15004 15264
rect 15068 15200 15084 15264
rect 15148 15200 15156 15264
rect 14836 14176 15156 15200
rect 14836 14112 14844 14176
rect 14908 14112 14924 14176
rect 14988 14112 15004 14176
rect 15068 14112 15084 14176
rect 15148 14112 15156 14176
rect 14836 13088 15156 14112
rect 14836 13024 14844 13088
rect 14908 13024 14924 13088
rect 14988 13024 15004 13088
rect 15068 13024 15084 13088
rect 15148 13024 15156 13088
rect 14836 12000 15156 13024
rect 14836 11936 14844 12000
rect 14908 11936 14924 12000
rect 14988 11936 15004 12000
rect 15068 11936 15084 12000
rect 15148 11936 15156 12000
rect 14836 10912 15156 11936
rect 14836 10848 14844 10912
rect 14908 10848 14924 10912
rect 14988 10848 15004 10912
rect 15068 10848 15084 10912
rect 15148 10848 15156 10912
rect 14836 9824 15156 10848
rect 14836 9760 14844 9824
rect 14908 9760 14924 9824
rect 14988 9760 15004 9824
rect 15068 9760 15084 9824
rect 15148 9760 15156 9824
rect 14836 8736 15156 9760
rect 14836 8672 14844 8736
rect 14908 8672 14924 8736
rect 14988 8672 15004 8736
rect 15068 8672 15084 8736
rect 15148 8672 15156 8736
rect 14836 7648 15156 8672
rect 14836 7584 14844 7648
rect 14908 7584 14924 7648
rect 14988 7584 15004 7648
rect 15068 7584 15084 7648
rect 15148 7584 15156 7648
rect 14836 6870 15156 7584
rect 14836 6634 14878 6870
rect 15114 6634 15156 6870
rect 14836 6560 15156 6634
rect 14836 6496 14844 6560
rect 14908 6496 14924 6560
rect 14988 6496 15004 6560
rect 15068 6496 15084 6560
rect 15148 6496 15156 6560
rect 14836 5472 15156 6496
rect 14836 5408 14844 5472
rect 14908 5408 14924 5472
rect 14988 5408 15004 5472
rect 15068 5408 15084 5472
rect 15148 5408 15156 5472
rect 14836 4384 15156 5408
rect 14836 4320 14844 4384
rect 14908 4320 14924 4384
rect 14988 4320 15004 4384
rect 15068 4320 15084 4384
rect 15148 4320 15156 4384
rect 14836 3296 15156 4320
rect 14836 3232 14844 3296
rect 14908 3232 14924 3296
rect 14988 3232 15004 3296
rect 15068 3232 15084 3296
rect 15148 3232 15156 3296
rect 14836 2208 15156 3232
rect 14836 2144 14844 2208
rect 14908 2144 14924 2208
rect 14988 2144 15004 2208
rect 15068 2144 15084 2208
rect 15148 2144 15156 2208
rect 14836 2128 15156 2144
rect 19466 29952 19787 29968
rect 19466 29888 19474 29952
rect 19538 29888 19554 29952
rect 19618 29888 19634 29952
rect 19698 29888 19714 29952
rect 19778 29888 19787 29952
rect 19466 28864 19787 29888
rect 19466 28800 19474 28864
rect 19538 28800 19554 28864
rect 19618 28800 19634 28864
rect 19698 28800 19714 28864
rect 19778 28800 19787 28864
rect 19466 27776 19787 28800
rect 19466 27712 19474 27776
rect 19538 27712 19554 27776
rect 19618 27712 19634 27776
rect 19698 27712 19714 27776
rect 19778 27712 19787 27776
rect 19466 26688 19787 27712
rect 19466 26624 19474 26688
rect 19538 26624 19554 26688
rect 19618 26624 19634 26688
rect 19698 26624 19714 26688
rect 19778 26624 19787 26688
rect 19466 25600 19787 26624
rect 19466 25536 19474 25600
rect 19538 25536 19554 25600
rect 19618 25536 19634 25600
rect 19698 25536 19714 25600
rect 19778 25536 19787 25600
rect 19466 24512 19787 25536
rect 19466 24448 19474 24512
rect 19538 24448 19554 24512
rect 19618 24448 19634 24512
rect 19698 24448 19714 24512
rect 19778 24448 19787 24512
rect 19466 23424 19787 24448
rect 19466 23360 19474 23424
rect 19538 23360 19554 23424
rect 19618 23360 19634 23424
rect 19698 23360 19714 23424
rect 19778 23360 19787 23424
rect 19466 22336 19787 23360
rect 19466 22272 19474 22336
rect 19538 22272 19554 22336
rect 19618 22272 19634 22336
rect 19698 22272 19714 22336
rect 19778 22272 19787 22336
rect 19466 21248 19787 22272
rect 19466 21184 19474 21248
rect 19538 21184 19554 21248
rect 19618 21184 19634 21248
rect 19698 21184 19714 21248
rect 19778 21184 19787 21248
rect 19466 20742 19787 21184
rect 19466 20506 19508 20742
rect 19744 20506 19787 20742
rect 19466 20160 19787 20506
rect 19466 20096 19474 20160
rect 19538 20096 19554 20160
rect 19618 20096 19634 20160
rect 19698 20096 19714 20160
rect 19778 20096 19787 20160
rect 19466 19072 19787 20096
rect 19466 19008 19474 19072
rect 19538 19008 19554 19072
rect 19618 19008 19634 19072
rect 19698 19008 19714 19072
rect 19778 19008 19787 19072
rect 19466 17984 19787 19008
rect 19466 17920 19474 17984
rect 19538 17920 19554 17984
rect 19618 17920 19634 17984
rect 19698 17920 19714 17984
rect 19778 17920 19787 17984
rect 19466 16896 19787 17920
rect 19466 16832 19474 16896
rect 19538 16832 19554 16896
rect 19618 16832 19634 16896
rect 19698 16832 19714 16896
rect 19778 16832 19787 16896
rect 19466 15808 19787 16832
rect 19466 15744 19474 15808
rect 19538 15744 19554 15808
rect 19618 15744 19634 15808
rect 19698 15744 19714 15808
rect 19778 15744 19787 15808
rect 19466 14720 19787 15744
rect 19466 14656 19474 14720
rect 19538 14656 19554 14720
rect 19618 14656 19634 14720
rect 19698 14656 19714 14720
rect 19778 14656 19787 14720
rect 19466 13632 19787 14656
rect 19466 13568 19474 13632
rect 19538 13568 19554 13632
rect 19618 13568 19634 13632
rect 19698 13568 19714 13632
rect 19778 13568 19787 13632
rect 19466 12544 19787 13568
rect 19466 12480 19474 12544
rect 19538 12480 19554 12544
rect 19618 12480 19634 12544
rect 19698 12480 19714 12544
rect 19778 12480 19787 12544
rect 19466 11494 19787 12480
rect 19466 11456 19508 11494
rect 19744 11456 19787 11494
rect 19466 11392 19474 11456
rect 19778 11392 19787 11456
rect 19466 11258 19508 11392
rect 19744 11258 19787 11392
rect 19466 10368 19787 11258
rect 19466 10304 19474 10368
rect 19538 10304 19554 10368
rect 19618 10304 19634 10368
rect 19698 10304 19714 10368
rect 19778 10304 19787 10368
rect 19466 9280 19787 10304
rect 19466 9216 19474 9280
rect 19538 9216 19554 9280
rect 19618 9216 19634 9280
rect 19698 9216 19714 9280
rect 19778 9216 19787 9280
rect 19466 8192 19787 9216
rect 19466 8128 19474 8192
rect 19538 8128 19554 8192
rect 19618 8128 19634 8192
rect 19698 8128 19714 8192
rect 19778 8128 19787 8192
rect 19466 7104 19787 8128
rect 19466 7040 19474 7104
rect 19538 7040 19554 7104
rect 19618 7040 19634 7104
rect 19698 7040 19714 7104
rect 19778 7040 19787 7104
rect 19466 6016 19787 7040
rect 19466 5952 19474 6016
rect 19538 5952 19554 6016
rect 19618 5952 19634 6016
rect 19698 5952 19714 6016
rect 19778 5952 19787 6016
rect 19466 4928 19787 5952
rect 19466 4864 19474 4928
rect 19538 4864 19554 4928
rect 19618 4864 19634 4928
rect 19698 4864 19714 4928
rect 19778 4864 19787 4928
rect 19466 3840 19787 4864
rect 19466 3776 19474 3840
rect 19538 3776 19554 3840
rect 19618 3776 19634 3840
rect 19698 3776 19714 3840
rect 19778 3776 19787 3840
rect 19466 2752 19787 3776
rect 19466 2688 19474 2752
rect 19538 2688 19554 2752
rect 19618 2688 19634 2752
rect 19698 2688 19714 2752
rect 19778 2688 19787 2752
rect 19466 2128 19787 2688
rect 24097 29408 24417 29968
rect 24097 29344 24105 29408
rect 24169 29344 24185 29408
rect 24249 29344 24265 29408
rect 24329 29344 24345 29408
rect 24409 29344 24417 29408
rect 24097 28320 24417 29344
rect 24097 28256 24105 28320
rect 24169 28256 24185 28320
rect 24249 28256 24265 28320
rect 24329 28256 24345 28320
rect 24409 28256 24417 28320
rect 24097 27232 24417 28256
rect 24097 27168 24105 27232
rect 24169 27168 24185 27232
rect 24249 27168 24265 27232
rect 24329 27168 24345 27232
rect 24409 27168 24417 27232
rect 24097 26144 24417 27168
rect 24097 26080 24105 26144
rect 24169 26080 24185 26144
rect 24249 26080 24265 26144
rect 24329 26080 24345 26144
rect 24409 26080 24417 26144
rect 24097 25366 24417 26080
rect 24097 25130 24139 25366
rect 24375 25130 24417 25366
rect 24097 25056 24417 25130
rect 24097 24992 24105 25056
rect 24169 24992 24185 25056
rect 24249 24992 24265 25056
rect 24329 24992 24345 25056
rect 24409 24992 24417 25056
rect 24097 23968 24417 24992
rect 24097 23904 24105 23968
rect 24169 23904 24185 23968
rect 24249 23904 24265 23968
rect 24329 23904 24345 23968
rect 24409 23904 24417 23968
rect 24097 22880 24417 23904
rect 24097 22816 24105 22880
rect 24169 22816 24185 22880
rect 24249 22816 24265 22880
rect 24329 22816 24345 22880
rect 24409 22816 24417 22880
rect 24097 21792 24417 22816
rect 24097 21728 24105 21792
rect 24169 21728 24185 21792
rect 24249 21728 24265 21792
rect 24329 21728 24345 21792
rect 24409 21728 24417 21792
rect 24097 20704 24417 21728
rect 24097 20640 24105 20704
rect 24169 20640 24185 20704
rect 24249 20640 24265 20704
rect 24329 20640 24345 20704
rect 24409 20640 24417 20704
rect 24097 19616 24417 20640
rect 24097 19552 24105 19616
rect 24169 19552 24185 19616
rect 24249 19552 24265 19616
rect 24329 19552 24345 19616
rect 24409 19552 24417 19616
rect 24097 18528 24417 19552
rect 24097 18464 24105 18528
rect 24169 18464 24185 18528
rect 24249 18464 24265 18528
rect 24329 18464 24345 18528
rect 24409 18464 24417 18528
rect 24097 17440 24417 18464
rect 24097 17376 24105 17440
rect 24169 17376 24185 17440
rect 24249 17376 24265 17440
rect 24329 17376 24345 17440
rect 24409 17376 24417 17440
rect 24097 16352 24417 17376
rect 24097 16288 24105 16352
rect 24169 16288 24185 16352
rect 24249 16288 24265 16352
rect 24329 16288 24345 16352
rect 24409 16288 24417 16352
rect 24097 16118 24417 16288
rect 24097 15882 24139 16118
rect 24375 15882 24417 16118
rect 24097 15264 24417 15882
rect 24097 15200 24105 15264
rect 24169 15200 24185 15264
rect 24249 15200 24265 15264
rect 24329 15200 24345 15264
rect 24409 15200 24417 15264
rect 24097 14176 24417 15200
rect 24097 14112 24105 14176
rect 24169 14112 24185 14176
rect 24249 14112 24265 14176
rect 24329 14112 24345 14176
rect 24409 14112 24417 14176
rect 24097 13088 24417 14112
rect 24097 13024 24105 13088
rect 24169 13024 24185 13088
rect 24249 13024 24265 13088
rect 24329 13024 24345 13088
rect 24409 13024 24417 13088
rect 24097 12000 24417 13024
rect 24097 11936 24105 12000
rect 24169 11936 24185 12000
rect 24249 11936 24265 12000
rect 24329 11936 24345 12000
rect 24409 11936 24417 12000
rect 24097 10912 24417 11936
rect 24097 10848 24105 10912
rect 24169 10848 24185 10912
rect 24249 10848 24265 10912
rect 24329 10848 24345 10912
rect 24409 10848 24417 10912
rect 24097 9824 24417 10848
rect 24097 9760 24105 9824
rect 24169 9760 24185 9824
rect 24249 9760 24265 9824
rect 24329 9760 24345 9824
rect 24409 9760 24417 9824
rect 24097 8736 24417 9760
rect 24097 8672 24105 8736
rect 24169 8672 24185 8736
rect 24249 8672 24265 8736
rect 24329 8672 24345 8736
rect 24409 8672 24417 8736
rect 24097 7648 24417 8672
rect 24097 7584 24105 7648
rect 24169 7584 24185 7648
rect 24249 7584 24265 7648
rect 24329 7584 24345 7648
rect 24409 7584 24417 7648
rect 24097 6870 24417 7584
rect 24097 6634 24139 6870
rect 24375 6634 24417 6870
rect 24097 6560 24417 6634
rect 24097 6496 24105 6560
rect 24169 6496 24185 6560
rect 24249 6496 24265 6560
rect 24329 6496 24345 6560
rect 24409 6496 24417 6560
rect 24097 5472 24417 6496
rect 24097 5408 24105 5472
rect 24169 5408 24185 5472
rect 24249 5408 24265 5472
rect 24329 5408 24345 5472
rect 24409 5408 24417 5472
rect 24097 4384 24417 5408
rect 24097 4320 24105 4384
rect 24169 4320 24185 4384
rect 24249 4320 24265 4384
rect 24329 4320 24345 4384
rect 24409 4320 24417 4384
rect 24097 3296 24417 4320
rect 24097 3232 24105 3296
rect 24169 3232 24185 3296
rect 24249 3232 24265 3296
rect 24329 3232 24345 3296
rect 24409 3232 24417 3296
rect 24097 2208 24417 3232
rect 24097 2144 24105 2208
rect 24169 2144 24185 2208
rect 24249 2144 24265 2208
rect 24329 2144 24345 2208
rect 24409 2144 24417 2208
rect 24097 2128 24417 2144
<< via4 >>
rect 5616 25130 5852 25366
rect 5616 15882 5852 16118
rect 5616 6634 5852 6870
rect 10247 20506 10483 20742
rect 10247 11456 10483 11494
rect 10247 11392 10277 11456
rect 10277 11392 10293 11456
rect 10293 11392 10357 11456
rect 10357 11392 10373 11456
rect 10373 11392 10437 11456
rect 10437 11392 10453 11456
rect 10453 11392 10483 11456
rect 10247 11258 10483 11392
rect 14878 25130 15114 25366
rect 14878 15882 15114 16118
rect 14878 6634 15114 6870
rect 19508 20506 19744 20742
rect 19508 11456 19744 11494
rect 19508 11392 19538 11456
rect 19538 11392 19554 11456
rect 19554 11392 19618 11456
rect 19618 11392 19634 11456
rect 19634 11392 19698 11456
rect 19698 11392 19714 11456
rect 19714 11392 19744 11456
rect 19508 11258 19744 11392
rect 24139 25130 24375 25366
rect 24139 15882 24375 16118
rect 24139 6634 24375 6870
<< metal5 >>
rect 1104 25366 28888 25408
rect 1104 25130 5616 25366
rect 5852 25130 14878 25366
rect 15114 25130 24139 25366
rect 24375 25130 28888 25366
rect 1104 25088 28888 25130
rect 1104 20742 28888 20784
rect 1104 20506 10247 20742
rect 10483 20506 19508 20742
rect 19744 20506 28888 20742
rect 1104 20464 28888 20506
rect 1104 16118 28888 16160
rect 1104 15882 5616 16118
rect 5852 15882 14878 16118
rect 15114 15882 24139 16118
rect 24375 15882 28888 16118
rect 1104 15840 28888 15882
rect 1104 11494 28888 11536
rect 1104 11258 10247 11494
rect 10483 11258 19508 11494
rect 19744 11258 28888 11494
rect 1104 11216 28888 11258
rect 1104 6870 28888 6912
rect 1104 6634 5616 6870
rect 5852 6634 14878 6870
rect 15114 6634 24139 6870
rect 24375 6634 28888 6870
rect 1104 6592 28888 6634
use sky130_fd_sc_hd__buf_1  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1620791022
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_6
timestamp 1620791022
transform 1 0 1656 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 2760 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1620791022
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1620791022
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1620791022
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1620791022
transform 1 0 3864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26
timestamp 1620791022
transform 1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1620791022
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1620791022
transform 1 0 6532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42
timestamp 1620791022
transform 1 0 4968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1620791022
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1620791022
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1620791022
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_70
timestamp 1620791022
transform 1 0 7544 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_71
timestamp 1620791022
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1620791022
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1620791022
transform 1 0 9752 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_100
timestamp 1620791022
transform 1 0 10304 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1620791022
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1620791022
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2ai_1  _135_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 12788 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_1_119 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 12052 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_117
timestamp 1620791022
transform 1 0 11868 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1620791022
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1620791022
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1620791022
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1620791022
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_106
timestamp 1620791022
transform 1 0 10856 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _126_
timestamp 1620791022
transform -1 0 14168 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _125_
timestamp 1620791022
transform -1 0 13524 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_131
timestamp 1620791022
transform 1 0 13156 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_142
timestamp 1620791022
transform 1 0 14168 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_129
timestamp 1620791022
transform 1 0 12972 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1620791022
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1620791022
transform 1 0 13524 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_127
timestamp 1620791022
transform 1 0 12788 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1620791022
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1620791022
transform 1 0 15272 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_158
timestamp 1620791022
transform 1 0 15640 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_146
timestamp 1620791022
transform 1 0 14536 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_166
timestamp 1620791022
transform 1 0 16376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_170
timestamp 1620791022
transform 1 0 16744 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1620791022
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1620791022
transform 1 0 16928 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1620791022
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_175
timestamp 1620791022
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1620791022
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1620791022
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1620791022
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 20056 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_196
timestamp 1620791022
transform 1 0 19136 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_202
timestamp 1620791022
transform 1 0 19688 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_206
timestamp 1620791022
transform 1 0 20056 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1620791022
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1620791022
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_204
timestamp 1620791022
transform 1 0 19872 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 20700 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_226 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 21896 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_212
timestamp 1620791022
transform 1 0 20608 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_229
timestamp 1620791022
transform 1 0 22172 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_216
timestamp 1620791022
transform 1 0 20976 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1620791022
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1620791022
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_218
timestamp 1620791022
transform 1 0 21160 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_241
timestamp 1620791022
transform 1 0 23276 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_245
timestamp 1620791022
transform 1 0 23644 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_233
timestamp 1620791022
transform 1 0 22540 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1620791022
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_265
timestamp 1620791022
transform 1 0 25484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_253
timestamp 1620791022
transform 1 0 24380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_262
timestamp 1620791022
transform 1 0 25208 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1620791022
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_257
timestamp 1620791022
transform 1 0 24748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_277
timestamp 1620791022
transform 1 0 26588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_274
timestamp 1620791022
transform 1 0 26312 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_286
timestamp 1620791022
transform 1 0 27416 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1620791022
transform 1 0 27416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1620791022
transform 1 0 27324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_282
timestamp 1620791022
transform 1 0 27048 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1620791022
transform -1 0 27416 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_291
timestamp 1620791022
transform 1 0 27876 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1620791022
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1620791022
transform 1 0 27784 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp 1620791022
transform 1 0 28060 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1620791022
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1620791022
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1620791022
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1620791022
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1620791022
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1620791022
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1620791022
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1620791022
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1620791022
transform 1 0 6072 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1620791022
transform 1 0 4968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1620791022
transform 1 0 7176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_78
timestamp 1620791022
transform 1 0 8280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 10580 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1620791022
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1620791022
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1620791022
transform 1 0 10212 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _174_
timestamp 1620791022
transform -1 0 13892 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_119
timestamp 1620791022
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1620791022
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_139
timestamp 1620791022
transform 1 0 13892 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1620791022
transform 1 0 14352 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 15088 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_161
timestamp 1620791022
transform 1 0 15916 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_185
timestamp 1620791022
transform 1 0 18124 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_173
timestamp 1620791022
transform 1 0 17020 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1620791022
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1620791022
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1620791022
transform 1 0 19228 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_225
timestamp 1620791022
transform 1 0 21804 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_213
timestamp 1620791022
transform 1 0 20700 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_237
timestamp 1620791022
transform 1 0 22908 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_249
timestamp 1620791022
transform 1 0 24012 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_270
timestamp 1620791022
transform 1 0 25944 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_258
timestamp 1620791022
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1620791022
transform 1 0 24748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_282
timestamp 1620791022
transform 1 0 27048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1620791022
transform 1 0 28520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1620791022
transform 1 0 28152 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1620791022
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1620791022
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1620791022
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1620791022
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1620791022
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1620791022
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1620791022
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1620791022
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1620791022
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1620791022
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1620791022
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1620791022
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__a31oi_1  _131_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 12144 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _142_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 11224 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_119
timestamp 1620791022
transform 1 0 12052 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_106
timestamp 1620791022
transform 1 0 10856 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1620791022
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp 1620791022
transform 1 0 12604 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_115
timestamp 1620791022
transform 1 0 11684 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_110
timestamp 1620791022
transform 1 0 11224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _173_
timestamp 1620791022
transform 1 0 12972 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_3_145
timestamp 1620791022
transform 1 0 14444 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _165_
timestamp 1620791022
transform 1 0 14996 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1620791022
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1620791022
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1620791022
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_167
timestamp 1620791022
transform 1 0 16468 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1620791022
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1620791022
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_229
timestamp 1620791022
transform 1 0 22172 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1620791022
transform 1 0 22080 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_220
timestamp 1620791022
transform 1 0 21344 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_241
timestamp 1620791022
transform 1 0 23276 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_265
timestamp 1620791022
transform 1 0 25484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_253
timestamp 1620791022
transform 1 0 24380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_286
timestamp 1620791022
transform 1 0 27416 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1620791022
transform 1 0 27324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_277
timestamp 1620791022
transform 1 0 26588 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_298
timestamp 1620791022
transform 1 0 28520 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1620791022
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1620791022
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1620791022
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1620791022
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1620791022
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1620791022
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1620791022
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1620791022
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1620791022
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1620791022
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1620791022
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _175_
timestamp 1620791022
transform 1 0 10488 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _158_
timestamp 1620791022
transform -1 0 10120 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1620791022
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_98
timestamp 1620791022
transform 1 0 10120 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_87
timestamp 1620791022
transform 1 0 9108 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 12880 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_118
timestamp 1620791022
transform 1 0 11960 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 13248 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1620791022
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_144
timestamp 1620791022
transform 1 0 14352 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_139
timestamp 1620791022
transform 1 0 13892 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp 1620791022
transform 1 0 12880 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _162_
timestamp 1620791022
transform 1 0 15824 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _157_
timestamp 1620791022
transform 1 0 14720 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_159
timestamp 1620791022
transform 1 0 15732 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_151
timestamp 1620791022
transform 1 0 14996 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_181
timestamp 1620791022
transform 1 0 17756 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_169
timestamp 1620791022
transform 1 0 16652 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_193
timestamp 1620791022
transform 1 0 18860 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_199
timestamp 1620791022
transform 1 0 19412 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_201
timestamp 1620791022
transform 1 0 19596 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1620791022
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_225
timestamp 1620791022
transform 1 0 21804 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_213
timestamp 1620791022
transform 1 0 20700 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_237
timestamp 1620791022
transform 1 0 22908 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_249
timestamp 1620791022
transform 1 0 24012 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_270
timestamp 1620791022
transform 1 0 25944 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_258
timestamp 1620791022
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1620791022
transform 1 0 24748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_282
timestamp 1620791022
transform 1 0 27048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp 1620791022
transform 1 0 28520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_294
timestamp 1620791022
transform 1 0 28152 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1620791022
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1620791022
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1620791022
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1620791022
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1620791022
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1620791022
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_51
timestamp 1620791022
transform 1 0 5796 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1620791022
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1620791022
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1620791022
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1620791022
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1620791022
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 12236 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _153_
timestamp 1620791022
transform -1 0 11224 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_115
timestamp 1620791022
transform 1 0 11684 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_106
timestamp 1620791022
transform 1 0 10856 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1620791022
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_110
timestamp 1620791022
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _143_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 13248 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _141_
timestamp 1620791022
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1620791022
transform 1 0 13892 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_128
timestamp 1620791022
transform 1 0 12880 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp 1620791022
transform -1 0 16008 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1620791022
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_146
timestamp 1620791022
transform 1 0 14536 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_162
timestamp 1620791022
transform 1 0 16008 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_170
timestamp 1620791022
transform 1 0 16744 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1620791022
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_172
timestamp 1620791022
transform 1 0 16928 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1620791022
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1620791022
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1620791022
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_229
timestamp 1620791022
transform 1 0 22172 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1620791022
transform 1 0 22080 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_220
timestamp 1620791022
transform 1 0 21344 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_241
timestamp 1620791022
transform 1 0 23276 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_265
timestamp 1620791022
transform 1 0 25484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_253
timestamp 1620791022
transform 1 0 24380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_286
timestamp 1620791022
transform 1 0 27416 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1620791022
transform 1 0 27324 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_277
timestamp 1620791022
transform 1 0 26588 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_298
timestamp 1620791022
transform 1 0 28520 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1620791022
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1620791022
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1620791022
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1620791022
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1620791022
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1620791022
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1620791022
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1620791022
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1620791022
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1620791022
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1620791022
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1620791022
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1620791022
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1620791022
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1620791022
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1620791022
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1620791022
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1620791022
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1620791022
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1620791022
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1620791022
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1620791022
transform -1 0 10396 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 10672 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_6_103
timestamp 1620791022
transform 1 0 10580 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1620791022
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1620791022
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_101
timestamp 1620791022
transform 1 0 10396 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_94
timestamp 1620791022
transform 1 0 9752 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1620791022
transform 1 0 10212 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _138_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 12788 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _139_
timestamp 1620791022
transform -1 0 12788 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _130_
timestamp 1620791022
transform 1 0 10764 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _129_
timestamp 1620791022
transform -1 0 11960 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1620791022
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_115
timestamp 1620791022
transform 1 0 11684 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_110
timestamp 1620791022
transform 1 0 11224 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_118
timestamp 1620791022
transform 1 0 11960 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_109
timestamp 1620791022
transform 1 0 11132 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_134
timestamp 1620791022
transform 1 0 13432 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_127
timestamp 1620791022
transform 1 0 12788 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_127
timestamp 1620791022
transform 1 0 12788 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_131
timestamp 1620791022
transform 1 0 13156 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1620791022
transform -1 0 13432 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _132_
timestamp 1620791022
transform 1 0 13248 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_6_144
timestamp 1620791022
transform 1 0 14352 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1620791022
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_137
timestamp 1620791022
transform 1 0 13708 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _166_
timestamp 1620791022
transform 1 0 13800 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp 1620791022
transform -1 0 14996 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_154
timestamp 1620791022
transform 1 0 15272 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_163
timestamp 1620791022
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_151
timestamp 1620791022
transform 1 0 14996 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_166
timestamp 1620791022
transform 1 0 16376 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_170
timestamp 1620791022
transform 1 0 16744 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1620791022
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1620791022
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_187
timestamp 1620791022
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_175
timestamp 1620791022
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1620791022
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_199
timestamp 1620791022
transform 1 0 19412 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1620791022
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1620791022
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1620791022
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1620791022
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_229
timestamp 1620791022
transform 1 0 22172 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_225
timestamp 1620791022
transform 1 0 21804 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_213
timestamp 1620791022
transform 1 0 20700 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1620791022
transform 1 0 22080 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_220
timestamp 1620791022
transform 1 0 21344 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_241
timestamp 1620791022
transform 1 0 23276 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_237
timestamp 1620791022
transform 1 0 22908 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_249
timestamp 1620791022
transform 1 0 24012 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_265
timestamp 1620791022
transform 1 0 25484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_253
timestamp 1620791022
transform 1 0 24380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_270
timestamp 1620791022
transform 1 0 25944 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_258
timestamp 1620791022
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1620791022
transform 1 0 24748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_286
timestamp 1620791022
transform 1 0 27416 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_282
timestamp 1620791022
transform 1 0 27048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1620791022
transform 1 0 27324 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_277
timestamp 1620791022
transform 1 0 26588 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_298
timestamp 1620791022
transform 1 0 28520 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1620791022
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_294
timestamp 1620791022
transform 1 0 28152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1620791022
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1620791022
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1620791022
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1620791022
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1620791022
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1620791022
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1620791022
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1620791022
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1620791022
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1620791022
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1620791022
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1620791022
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _167_
timestamp 1620791022
transform -1 0 11776 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1620791022
transform 1 0 10212 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1620791022
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1620791022
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 12236 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_120
timestamp 1620791022
transform 1 0 12144 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_116
timestamp 1620791022
transform 1 0 11776 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 13432 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1620791022
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_144
timestamp 1620791022
transform 1 0 14352 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_139
timestamp 1620791022
transform 1 0 13892 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_130
timestamp 1620791022
transform 1 0 13064 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _137_
timestamp 1620791022
transform 1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _112_
timestamp 1620791022
transform -1 0 14996 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_158
timestamp 1620791022
transform 1 0 15640 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_151
timestamp 1620791022
transform 1 0 14996 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_182
timestamp 1620791022
transform 1 0 17848 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_170
timestamp 1620791022
transform 1 0 16744 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_194
timestamp 1620791022
transform 1 0 18952 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1620791022
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1620791022
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_225
timestamp 1620791022
transform 1 0 21804 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_213
timestamp 1620791022
transform 1 0 20700 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_237
timestamp 1620791022
transform 1 0 22908 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_249
timestamp 1620791022
transform 1 0 24012 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_270
timestamp 1620791022
transform 1 0 25944 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_258
timestamp 1620791022
transform 1 0 24840 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1620791022
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_282
timestamp 1620791022
transform 1 0 27048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1620791022
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_294
timestamp 1620791022
transform 1 0 28152 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1620791022
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1620791022
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1620791022
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1620791022
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1620791022
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1620791022
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51
timestamp 1620791022
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1620791022
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1620791022
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1620791022
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1620791022
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _168_
timestamp 1620791022
transform -1 0 11224 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__and3_1  _133_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 12052 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1620791022
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_115
timestamp 1620791022
transform 1 0 11684 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_110
timestamp 1620791022
transform 1 0 11224 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_124
timestamp 1620791022
transform 1 0 12512 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _100_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 14812 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_132
timestamp 1620791022
transform 1 0 13248 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _090_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 13708 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_137
timestamp 1620791022
transform 1 0 13708 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 15180 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_156
timestamp 1620791022
transform 1 0 15456 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_149
timestamp 1620791022
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1620791022
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1620791022
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1620791022
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_168
timestamp 1620791022
transform 1 0 16560 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1620791022
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1620791022
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_229
timestamp 1620791022
transform 1 0 22172 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1620791022
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_220
timestamp 1620791022
transform 1 0 21344 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_241
timestamp 1620791022
transform 1 0 23276 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_265
timestamp 1620791022
transform 1 0 25484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_253
timestamp 1620791022
transform 1 0 24380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_286
timestamp 1620791022
transform 1 0 27416 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1620791022
transform 1 0 27324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_277
timestamp 1620791022
transform 1 0 26588 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_298
timestamp 1620791022
transform 1 0 28520 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1620791022
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1620791022
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1620791022
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1620791022
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1620791022
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1620791022
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1620791022
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1620791022
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1620791022
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1620791022
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1620791022
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 10580 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_10_87
timestamp 1620791022
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1620791022
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_99
timestamp 1620791022
transform 1 0 10212 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _144_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 12880 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _134_
timestamp 1620791022
transform 1 0 11684 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_10_108
timestamp 1620791022
transform 1 0 11040 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_114
timestamp 1620791022
transform 1 0 11592 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_120
timestamp 1620791022
transform 1 0 12144 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _101_
timestamp 1620791022
transform -1 0 13524 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1620791022
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1620791022
transform 1 0 14352 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1620791022
transform 1 0 12880 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1620791022
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _177_
timestamp 1620791022
transform 1 0 14720 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_10_164
timestamp 1620791022
transform 1 0 16192 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_176
timestamp 1620791022
transform 1 0 17296 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1620791022
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_188
timestamp 1620791022
transform 1 0 18400 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1620791022
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_225
timestamp 1620791022
transform 1 0 21804 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_213
timestamp 1620791022
transform 1 0 20700 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_237
timestamp 1620791022
transform 1 0 22908 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_249
timestamp 1620791022
transform 1 0 24012 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_270
timestamp 1620791022
transform 1 0 25944 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_258
timestamp 1620791022
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1620791022
transform 1 0 24748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_282
timestamp 1620791022
transform 1 0 27048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1620791022
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_294
timestamp 1620791022
transform 1 0 28152 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1620791022
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1620791022
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1620791022
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1620791022
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1620791022
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1620791022
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1620791022
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1620791022
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1620791022
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_82
timestamp 1620791022
transform 1 0 8648 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1620791022
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_94
timestamp 1620791022
transform 1 0 9752 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_102
timestamp 1620791022
transform 1 0 10488 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _107_
timestamp 1620791022
transform -1 0 12328 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _151_
timestamp 1620791022
transform -1 0 11040 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_108
timestamp 1620791022
transform 1 0 11040 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_122
timestamp 1620791022
transform 1 0 12328 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1620791022
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1620791022
transform 1 0 11684 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1620791022
transform -1 0 13892 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_134
timestamp 1620791022
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_139
timestamp 1620791022
transform 1 0 13892 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_145
timestamp 1620791022
transform 1 0 14444 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _094_
timestamp 1620791022
transform 1 0 15180 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _093_
timestamp 1620791022
transform 1 0 14536 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_156
timestamp 1620791022
transform 1 0 15456 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_149
timestamp 1620791022
transform 1 0 14812 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1620791022
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1620791022
transform 1 0 16928 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1620791022
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_168
timestamp 1620791022
transform 1 0 16560 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1620791022
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1620791022
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_229
timestamp 1620791022
transform 1 0 22172 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1620791022
transform 1 0 22080 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_220
timestamp 1620791022
transform 1 0 21344 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_241
timestamp 1620791022
transform 1 0 23276 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_265
timestamp 1620791022
transform 1 0 25484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_253
timestamp 1620791022
transform 1 0 24380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_286
timestamp 1620791022
transform 1 0 27416 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1620791022
transform 1 0 27324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_277
timestamp 1620791022
transform 1 0 26588 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_298
timestamp 1620791022
transform 1 0 28520 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1620791022
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1620791022
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1620791022
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1620791022
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1620791022
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1620791022
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1620791022
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1620791022
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1620791022
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_66
timestamp 1620791022
transform 1 0 7176 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_78
timestamp 1620791022
transform 1 0 8280 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _149_
timestamp 1620791022
transform -1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_99
timestamp 1620791022
transform 1 0 10212 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_87
timestamp 1620791022
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1620791022
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_103
timestamp 1620791022
transform 1 0 10580 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 10948 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 12052 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_12_115
timestamp 1620791022
transform 1 0 11684 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1620791022
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_144
timestamp 1620791022
transform 1 0 14352 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_139
timestamp 1620791022
transform 1 0 13892 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _178_
timestamp 1620791022
transform 1 0 14720 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_12_164
timestamp 1620791022
transform 1 0 16192 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_176
timestamp 1620791022
transform 1 0 17296 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1620791022
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_188
timestamp 1620791022
transform 1 0 18400 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1620791022
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_225
timestamp 1620791022
transform 1 0 21804 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_213
timestamp 1620791022
transform 1 0 20700 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_237
timestamp 1620791022
transform 1 0 22908 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_249
timestamp 1620791022
transform 1 0 24012 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_270
timestamp 1620791022
transform 1 0 25944 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_258
timestamp 1620791022
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1620791022
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_282
timestamp 1620791022
transform 1 0 27048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp 1620791022
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_294
timestamp 1620791022
transform 1 0 28152 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1620791022
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1620791022
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1620791022
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1620791022
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1620791022
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1620791022
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1620791022
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1620791022
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1620791022
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1620791022
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1620791022
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1620791022
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_51
timestamp 1620791022
transform 1 0 5796 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1620791022
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1620791022
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1620791022
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1620791022
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1620791022
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1620791022
transform 1 0 8648 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1620791022
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_78
timestamp 1620791022
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _180_
timestamp 1620791022
transform 1 0 10028 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _179_
timestamp 1620791022
transform 1 0 9752 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_95
timestamp 1620791022
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1620791022
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_87
timestamp 1620791022
transform 1 0 9108 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 12420 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _113_
timestamp 1620791022
transform -1 0 12328 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1620791022
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1620791022
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_122
timestamp 1620791022
transform 1 0 12328 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_113
timestamp 1620791022
transform 1 0 11500 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1620791022
transform 1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_110
timestamp 1620791022
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _116_
timestamp 1620791022
transform 1 0 12696 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_13_135
timestamp 1620791022
transform 1 0 13524 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_131
timestamp 1620791022
transform 1 0 13156 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_135
timestamp 1620791022
transform 1 0 13524 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1620791022
transform -1 0 13892 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_139
timestamp 1620791022
transform 1 0 13892 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_141
timestamp 1620791022
transform 1 0 14076 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _104_
timestamp 1620791022
transform 1 0 13800 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_144
timestamp 1620791022
transform 1 0 14352 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1620791022
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _096_
timestamp 1620791022
transform -1 0 14904 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _095_
timestamp 1620791022
transform -1 0 15640 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _170_
timestamp 1620791022
transform 1 0 14720 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _159_
timestamp 1620791022
transform 1 0 16008 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_165
timestamp 1620791022
transform 1 0 16284 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_164
timestamp 1620791022
transform 1 0 16192 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_158
timestamp 1620791022
transform 1 0 15640 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_150
timestamp 1620791022
transform 1 0 14904 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_176
timestamp 1620791022
transform 1 0 17296 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1620791022
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1620791022
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1620791022
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1620791022
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_188
timestamp 1620791022
transform 1 0 18400 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1620791022
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1620791022
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1620791022
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_225
timestamp 1620791022
transform 1 0 21804 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_213
timestamp 1620791022
transform 1 0 20700 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_229
timestamp 1620791022
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1620791022
transform 1 0 22080 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_220
timestamp 1620791022
transform 1 0 21344 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_237
timestamp 1620791022
transform 1 0 22908 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_241
timestamp 1620791022
transform 1 0 23276 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_249
timestamp 1620791022
transform 1 0 24012 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_270
timestamp 1620791022
transform 1 0 25944 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_258
timestamp 1620791022
transform 1 0 24840 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_265
timestamp 1620791022
transform 1 0 25484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_253
timestamp 1620791022
transform 1 0 24380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1620791022
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_282
timestamp 1620791022
transform 1 0 27048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_286
timestamp 1620791022
transform 1 0 27416 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1620791022
transform 1 0 27324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_277
timestamp 1620791022
transform 1 0 26588 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_298
timestamp 1620791022
transform 1 0 28520 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_298
timestamp 1620791022
transform 1 0 28520 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_294
timestamp 1620791022
transform 1 0 28152 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1620791022
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1620791022
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1620791022
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1620791022
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1620791022
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1620791022
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1620791022
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1620791022
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1620791022
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1620791022
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_82
timestamp 1620791022
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1620791022
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _117_
timestamp 1620791022
transform -1 0 10396 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_15_94
timestamp 1620791022
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_101
timestamp 1620791022
transform 1 0 10396 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 12880 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _111_
timestamp 1620791022
transform 1 0 10764 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1620791022
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1620791022
transform 1 0 11684 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_110
timestamp 1620791022
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_2  _124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 13892 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _097_
timestamp 1620791022
transform -1 0 13524 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_135
timestamp 1620791022
transform 1 0 13524 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_128
timestamp 1620791022
transform 1 0 12880 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _105_
timestamp 1620791022
transform -1 0 16192 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _102_
timestamp 1620791022
transform -1 0 15364 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_15_164
timestamp 1620791022
transform 1 0 16192 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_155
timestamp 1620791022
transform 1 0 15364 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_146
timestamp 1620791022
transform 1 0 14536 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_170
timestamp 1620791022
transform 1 0 16744 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1620791022
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1620791022
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1620791022
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1620791022
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1620791022
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_229
timestamp 1620791022
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1620791022
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_220
timestamp 1620791022
transform 1 0 21344 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_241
timestamp 1620791022
transform 1 0 23276 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_265
timestamp 1620791022
transform 1 0 25484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_253
timestamp 1620791022
transform 1 0 24380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_286
timestamp 1620791022
transform 1 0 27416 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1620791022
transform 1 0 27324 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_277
timestamp 1620791022
transform 1 0 26588 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_298
timestamp 1620791022
transform 1 0 28520 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1620791022
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1620791022
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1620791022
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1620791022
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1620791022
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1620791022
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1620791022
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_54
timestamp 1620791022
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1620791022
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_66
timestamp 1620791022
transform 1 0 7176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1620791022
transform 1 0 8280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _172_
timestamp 1620791022
transform -1 0 11132 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_16_87
timestamp 1620791022
transform 1 0 9108 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1620791022
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _109_
timestamp 1620791022
transform -1 0 11960 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _114_
timestamp 1620791022
transform 1 0 12328 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp 1620791022
transform 1 0 11960 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1620791022
transform 1 0 11132 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _120_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform 1 0 13340 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_127
timestamp 1620791022
transform 1 0 12788 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1620791022
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_144
timestamp 1620791022
transform 1 0 14352 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_139
timestamp 1620791022
transform 1 0 13892 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _169_
timestamp 1620791022
transform 1 0 14720 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_16_164
timestamp 1620791022
transform 1 0 16192 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_176
timestamp 1620791022
transform 1 0 17296 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1620791022
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_188
timestamp 1620791022
transform 1 0 18400 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1620791022
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_225
timestamp 1620791022
transform 1 0 21804 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_213
timestamp 1620791022
transform 1 0 20700 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_237
timestamp 1620791022
transform 1 0 22908 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_249
timestamp 1620791022
transform 1 0 24012 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_270
timestamp 1620791022
transform 1 0 25944 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_258
timestamp 1620791022
transform 1 0 24840 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1620791022
transform 1 0 24748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_282
timestamp 1620791022
transform 1 0 27048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_298
timestamp 1620791022
transform 1 0 28520 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_294
timestamp 1620791022
transform 1 0 28152 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1620791022
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1620791022
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1620791022
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1620791022
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1620791022
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1620791022
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1620791022
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1620791022
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1620791022
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_70
timestamp 1620791022
transform 1 0 7544 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_82
timestamp 1620791022
transform 1 0 8648 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _150_
timestamp 1620791022
transform 1 0 10304 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1620791022
transform -1 0 9936 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_96
timestamp 1620791022
transform 1 0 9936 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_90
timestamp 1620791022
transform 1 0 9384 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _121_
timestamp 1620791022
transform 1 0 12052 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1620791022
transform 1 0 11500 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1620791022
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1620791022
transform 1 0 11684 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_105
timestamp 1620791022
transform 1 0 10764 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _123_
timestamp 1620791022
transform 1 0 14260 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _146_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 13708 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_17_137
timestamp 1620791022
transform 1 0 13708 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_128
timestamp 1620791022
transform 1 0 12880 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _098_
timestamp 1620791022
transform -1 0 15732 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1620791022
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_152
timestamp 1620791022
transform 1 0 15088 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1620791022
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1620791022
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1620791022
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1620791022
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1620791022
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_229
timestamp 1620791022
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1620791022
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_220
timestamp 1620791022
transform 1 0 21344 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_241
timestamp 1620791022
transform 1 0 23276 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_265
timestamp 1620791022
transform 1 0 25484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_253
timestamp 1620791022
transform 1 0 24380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_286
timestamp 1620791022
transform 1 0 27416 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1620791022
transform 1 0 27324 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_277
timestamp 1620791022
transform 1 0 26588 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_298
timestamp 1620791022
transform 1 0 28520 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1620791022
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1620791022
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1620791022
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1620791022
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1620791022
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1620791022
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1620791022
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_54
timestamp 1620791022
transform 1 0 6072 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1620791022
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_66
timestamp 1620791022
transform 1 0 7176 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_78
timestamp 1620791022
transform 1 0 8280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _171_
timestamp 1620791022
transform 1 0 10212 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1620791022
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1620791022
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _148_
timestamp 1620791022
transform 1 0 12604 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_18_123
timestamp 1620791022
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_115
timestamp 1620791022
transform 1 0 11684 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1620791022
transform -1 0 13892 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1620791022
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_144
timestamp 1620791022
transform 1 0 14352 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_139
timestamp 1620791022
transform 1 0 13892 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_132
timestamp 1620791022
transform 1 0 13248 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _122_
timestamp 1620791022
transform -1 0 14996 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_163
timestamp 1620791022
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_151
timestamp 1620791022
transform 1 0 14996 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_187
timestamp 1620791022
transform 1 0 18308 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_175
timestamp 1620791022
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_199
timestamp 1620791022
transform 1 0 19412 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_201
timestamp 1620791022
transform 1 0 19596 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1620791022
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_225
timestamp 1620791022
transform 1 0 21804 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_213
timestamp 1620791022
transform 1 0 20700 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_237
timestamp 1620791022
transform 1 0 22908 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_249
timestamp 1620791022
transform 1 0 24012 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_270
timestamp 1620791022
transform 1 0 25944 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_258
timestamp 1620791022
transform 1 0 24840 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1620791022
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_282
timestamp 1620791022
transform 1 0 27048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_298
timestamp 1620791022
transform 1 0 28520 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_294
timestamp 1620791022
transform 1 0 28152 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1620791022
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1620791022
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1620791022
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1620791022
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1620791022
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1620791022
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1620791022
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1620791022
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1620791022
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1620791022
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1620791022
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1620791022
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1620791022
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_54
timestamp 1620791022
transform 1 0 6072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1620791022
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1620791022
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1620791022
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_66
timestamp 1620791022
transform 1 0 7176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1620791022
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1620791022
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_78
timestamp 1620791022
transform 1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_99
timestamp 1620791022
transform 1 0 10212 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1620791022
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1620791022
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1620791022
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_110
timestamp 1620791022
transform 1 0 11224 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1620791022
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_114
timestamp 1620791022
transform 1 0 11592 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_106
timestamp 1620791022
transform 1 0 10856 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_108
timestamp 1620791022
transform 1 0 11040 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1620791022
transform 1 0 10948 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _084_
timestamp 1620791022
transform 1 0 10764 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_122
timestamp 1620791022
transform 1 0 12328 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_115
timestamp 1620791022
transform 1 0 11684 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1620791022
transform 1 0 12052 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a31o_1  _085_
timestamp 1620791022
transform 1 0 11684 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _181_
timestamp 1620791022
transform 1 0 12144 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__o21a_1  _160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1620791022
transform -1 0 13708 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _161_
timestamp 1620791022
transform 1 0 13984 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_20_137
timestamp 1620791022
transform 1 0 13708 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_130
timestamp 1620791022
transform 1 0 13064 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1620791022
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_145
timestamp 1620791022
transform 1 0 14444 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1620791022
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_136
timestamp 1620791022
transform 1 0 13616 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1620791022
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_157
timestamp 1620791022
transform 1 0 15548 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1620791022
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_180
timestamp 1620791022
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_168
timestamp 1620791022
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1620791022
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1620791022
transform 1 0 16928 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1620791022
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1620791022
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1620791022
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1620791022
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1620791022
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_192
timestamp 1620791022
transform 1 0 18768 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_225
timestamp 1620791022
transform 1 0 21804 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_213
timestamp 1620791022
transform 1 0 20700 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_229
timestamp 1620791022
transform 1 0 22172 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1620791022
transform 1 0 22080 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_220
timestamp 1620791022
transform 1 0 21344 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_237
timestamp 1620791022
transform 1 0 22908 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_241
timestamp 1620791022
transform 1 0 23276 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_249
timestamp 1620791022
transform 1 0 24012 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_270
timestamp 1620791022
transform 1 0 25944 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_258
timestamp 1620791022
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_265
timestamp 1620791022
transform 1 0 25484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_253
timestamp 1620791022
transform 1 0 24380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1620791022
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_282
timestamp 1620791022
transform 1 0 27048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_286
timestamp 1620791022
transform 1 0 27416 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1620791022
transform 1 0 27324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_277
timestamp 1620791022
transform 1 0 26588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_298
timestamp 1620791022
transform 1 0 28520 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_298
timestamp 1620791022
transform 1 0 28520 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_294
timestamp 1620791022
transform 1 0 28152 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1620791022
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1620791022
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1620791022
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1620791022
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1620791022
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1620791022
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1620791022
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1620791022
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1620791022
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1620791022
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1620791022
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1620791022
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1620791022
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _147_
timestamp 1620791022
transform -1 0 11224 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _164_
timestamp 1620791022
transform -1 0 13524 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_106
timestamp 1620791022
transform 1 0 10856 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1620791022
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_115
timestamp 1620791022
transform 1 0 11684 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_110
timestamp 1620791022
transform 1 0 11224 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _182_
timestamp 1620791022
transform 1 0 13892 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_135
timestamp 1620791022
transform 1 0 13524 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_155
timestamp 1620791022
transform 1 0 15364 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1620791022
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_172
timestamp 1620791022
transform 1 0 16928 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1620791022
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_167
timestamp 1620791022
transform 1 0 16468 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1620791022
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1620791022
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_229
timestamp 1620791022
transform 1 0 22172 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1620791022
transform 1 0 22080 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_220
timestamp 1620791022
transform 1 0 21344 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_241
timestamp 1620791022
transform 1 0 23276 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_265
timestamp 1620791022
transform 1 0 25484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_253
timestamp 1620791022
transform 1 0 24380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_286
timestamp 1620791022
transform 1 0 27416 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1620791022
transform 1 0 27324 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_277
timestamp 1620791022
transform 1 0 26588 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_298
timestamp 1620791022
transform 1 0 28520 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1620791022
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1620791022
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1620791022
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1620791022
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1620791022
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1620791022
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1620791022
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1620791022
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1620791022
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_66
timestamp 1620791022
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1620791022
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1620791022
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1620791022
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1620791022
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _086_
timestamp 1620791022
transform -1 0 13340 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _083_
timestamp 1620791022
transform -1 0 12236 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_111
timestamp 1620791022
transform 1 0 11316 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_117
timestamp 1620791022
transform 1 0 11868 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_121
timestamp 1620791022
transform 1 0 12236 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1620791022
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1620791022
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1620791022
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_133
timestamp 1620791022
transform 1 0 13340 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1620791022
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_180
timestamp 1620791022
transform 1 0 17664 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1620791022
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1620791022
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1620791022
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_192
timestamp 1620791022
transform 1 0 18768 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_225
timestamp 1620791022
transform 1 0 21804 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_213
timestamp 1620791022
transform 1 0 20700 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_237
timestamp 1620791022
transform 1 0 22908 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_249
timestamp 1620791022
transform 1 0 24012 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_270
timestamp 1620791022
transform 1 0 25944 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_258
timestamp 1620791022
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1620791022
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_282
timestamp 1620791022
transform 1 0 27048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_298
timestamp 1620791022
transform 1 0 28520 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_294
timestamp 1620791022
transform 1 0 28152 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1620791022
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1620791022
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_18
timestamp 1620791022
transform 1 0 2760 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_6
timestamp 1620791022
transform 1 0 1656 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1620791022
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_30
timestamp 1620791022
transform 1 0 3864 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_58
timestamp 1620791022
transform 1 0 6440 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_42
timestamp 1620791022
transform 1 0 4968 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1620791022
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_54
timestamp 1620791022
transform 1 0 6072 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_82
timestamp 1620791022
transform 1 0 8648 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_70
timestamp 1620791022
transform 1 0 7544 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_94
timestamp 1620791022
transform 1 0 9752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _087_
timestamp 1620791022
transform -1 0 12420 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1620791022
transform 1 0 12052 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1620791022
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_123
timestamp 1620791022
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_115
timestamp 1620791022
transform 1 0 11684 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1620791022
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _088_
timestamp 1620791022
transform -1 0 13524 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1620791022
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1620791022
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1620791022
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1620791022
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1620791022
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1620791022
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1620791022
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1620791022
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_229
timestamp 1620791022
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1620791022
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_220
timestamp 1620791022
transform 1 0 21344 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_241
timestamp 1620791022
transform 1 0 23276 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_265
timestamp 1620791022
transform 1 0 25484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_253
timestamp 1620791022
transform 1 0 24380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_286
timestamp 1620791022
transform 1 0 27416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1620791022
transform 1 0 27324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_277
timestamp 1620791022
transform 1 0 26588 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_298
timestamp 1620791022
transform 1 0 28520 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1620791022
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1620791022
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1620791022
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1620791022
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1620791022
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1620791022
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1620791022
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1620791022
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1620791022
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1620791022
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_78
timestamp 1620791022
transform 1 0 8280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1620791022
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1620791022
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1620791022
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1620791022
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1620791022
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1620791022
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 1620791022
transform 1 0 14352 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1620791022
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _082_
timestamp 1620791022
transform -1 0 14996 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_163
timestamp 1620791022
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_151
timestamp 1620791022
transform 1 0 14996 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_187
timestamp 1620791022
transform 1 0 18308 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_175
timestamp 1620791022
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_199
timestamp 1620791022
transform 1 0 19412 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1620791022
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1620791022
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_225
timestamp 1620791022
transform 1 0 21804 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_213
timestamp 1620791022
transform 1 0 20700 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_237
timestamp 1620791022
transform 1 0 22908 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_249
timestamp 1620791022
transform 1 0 24012 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_270
timestamp 1620791022
transform 1 0 25944 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_258
timestamp 1620791022
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1620791022
transform 1 0 24748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_282
timestamp 1620791022
transform 1 0 27048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_298
timestamp 1620791022
transform 1 0 28520 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_294
timestamp 1620791022
transform 1 0 28152 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1620791022
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1620791022
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1620791022
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1620791022
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1620791022
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1620791022
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_51
timestamp 1620791022
transform 1 0 5796 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_58
timestamp 1620791022
transform 1 0 6440 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1620791022
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_82
timestamp 1620791022
transform 1 0 8648 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_70
timestamp 1620791022
transform 1 0 7544 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_94
timestamp 1620791022
transform 1 0 9752 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1620791022
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1620791022
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_106
timestamp 1620791022
transform 1 0 10856 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_139
timestamp 1620791022
transform 1 0 13892 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1620791022
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_151
timestamp 1620791022
transform 1 0 14996 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_163
timestamp 1620791022
transform 1 0 16100 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1620791022
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1620791022
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1620791022
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1620791022
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1620791022
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_229
timestamp 1620791022
transform 1 0 22172 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1620791022
transform 1 0 22080 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_220
timestamp 1620791022
transform 1 0 21344 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_241
timestamp 1620791022
transform 1 0 23276 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_265
timestamp 1620791022
transform 1 0 25484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_253
timestamp 1620791022
transform 1 0 24380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_286
timestamp 1620791022
transform 1 0 27416 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1620791022
transform 1 0 27324 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_277
timestamp 1620791022
transform 1 0 26588 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_298
timestamp 1620791022
transform 1 0 28520 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1620791022
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1620791022
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1620791022
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1620791022
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1620791022
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1620791022
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1620791022
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1620791022
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1620791022
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1620791022
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1620791022
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1620791022
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_51
timestamp 1620791022
transform 1 0 5796 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_58
timestamp 1620791022
transform 1 0 6440 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1620791022
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1620791022
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1620791022
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_82
timestamp 1620791022
transform 1 0 8648 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_70
timestamp 1620791022
transform 1 0 7544 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1620791022
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1620791022
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1620791022
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1620791022
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1620791022
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1620791022
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_115
timestamp 1620791022
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1620791022
transform 1 0 12420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_111
timestamp 1620791022
transform 1 0 11316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1620791022
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_106
timestamp 1620791022
transform 1 0 10856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_139
timestamp 1620791022
transform 1 0 13892 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_127
timestamp 1620791022
transform 1 0 12788 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1620791022
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1620791022
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1620791022
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_151
timestamp 1620791022
transform 1 0 14996 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1620791022
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_163
timestamp 1620791022
transform 1 0 16100 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1620791022
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1620791022
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_180
timestamp 1620791022
transform 1 0 17664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1620791022
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1620791022
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1620791022
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1620791022
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_201
timestamp 1620791022
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1620791022
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_192
timestamp 1620791022
transform 1 0 18768 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_229
timestamp 1620791022
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_225
timestamp 1620791022
transform 1 0 21804 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_213
timestamp 1620791022
transform 1 0 20700 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1620791022
transform 1 0 22080 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_220
timestamp 1620791022
transform 1 0 21344 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_241
timestamp 1620791022
transform 1 0 23276 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_237
timestamp 1620791022
transform 1 0 22908 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_249
timestamp 1620791022
transform 1 0 24012 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_265
timestamp 1620791022
transform 1 0 25484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_253
timestamp 1620791022
transform 1 0 24380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_270
timestamp 1620791022
transform 1 0 25944 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_258
timestamp 1620791022
transform 1 0 24840 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1620791022
transform 1 0 24748 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_290
timestamp 1620791022
transform 1 0 27784 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_282
timestamp 1620791022
transform 1 0 27048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1620791022
transform 1 0 27324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output9
timestamp 1620791022
transform 1 0 27876 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1620791022
transform 1 0 27416 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_277
timestamp 1620791022
transform 1 0 26588 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_298
timestamp 1620791022
transform 1 0 28520 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_295
timestamp 1620791022
transform 1 0 28244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_294
timestamp 1620791022
transform 1 0 28152 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1620791022
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1620791022
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1620791022
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1620791022
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1620791022
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1620791022
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1620791022
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1620791022
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_54
timestamp 1620791022
transform 1 0 6072 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1620791022
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1620791022
transform 1 0 7176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_78
timestamp 1620791022
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_99
timestamp 1620791022
transform 1 0 10212 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_87
timestamp 1620791022
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1620791022
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1620791022
transform 1 0 12420 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_111
timestamp 1620791022
transform 1 0 11316 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1620791022
transform 1 0 14352 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1620791022
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_135
timestamp 1620791022
transform 1 0 13524 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1620791022
transform 1 0 15456 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1620791022
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1620791022
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1620791022
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1620791022
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_192
timestamp 1620791022
transform 1 0 18768 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_225
timestamp 1620791022
transform 1 0 21804 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_213
timestamp 1620791022
transform 1 0 20700 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_237
timestamp 1620791022
transform 1 0 22908 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_249
timestamp 1620791022
transform 1 0 24012 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_270
timestamp 1620791022
transform 1 0 25944 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_258
timestamp 1620791022
transform 1 0 24840 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1620791022
transform 1 0 24748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_282
timestamp 1620791022
transform 1 0 27048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_298
timestamp 1620791022
transform 1 0 28520 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_294
timestamp 1620791022
transform 1 0 28152 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1620791022
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1620791022
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1620791022
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1620791022
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1620791022
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1620791022
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_51
timestamp 1620791022
transform 1 0 5796 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1620791022
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1620791022
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1620791022
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1620791022
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1620791022
transform 1 0 9752 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_115
timestamp 1620791022
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1620791022
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_106
timestamp 1620791022
transform 1 0 10856 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_139
timestamp 1620791022
transform 1 0 13892 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_127
timestamp 1620791022
transform 1 0 12788 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1620791022
transform 1 0 14996 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_163
timestamp 1620791022
transform 1 0 16100 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1620791022
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1620791022
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1620791022
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1620791022
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1620791022
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_229
timestamp 1620791022
transform 1 0 22172 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1620791022
transform 1 0 22080 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_220
timestamp 1620791022
transform 1 0 21344 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_241
timestamp 1620791022
transform 1 0 23276 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_265
timestamp 1620791022
transform 1 0 25484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_253
timestamp 1620791022
transform 1 0 24380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_286
timestamp 1620791022
transform 1 0 27416 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1620791022
transform 1 0 27324 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_277
timestamp 1620791022
transform 1 0 26588 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_298
timestamp 1620791022
transform 1 0 28520 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1620791022
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1620791022
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1620791022
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1620791022
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1620791022
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1620791022
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1620791022
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_54
timestamp 1620791022
transform 1 0 6072 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_42
timestamp 1620791022
transform 1 0 4968 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_66
timestamp 1620791022
transform 1 0 7176 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_78
timestamp 1620791022
transform 1 0 8280 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_99
timestamp 1620791022
transform 1 0 10212 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_87
timestamp 1620791022
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1620791022
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_123
timestamp 1620791022
transform 1 0 12420 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_111
timestamp 1620791022
transform 1 0 11316 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1620791022
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1620791022
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_135
timestamp 1620791022
transform 1 0 13524 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_156
timestamp 1620791022
transform 1 0 15456 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_180
timestamp 1620791022
transform 1 0 17664 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1620791022
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1620791022
transform 1 0 19596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1620791022
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_192
timestamp 1620791022
transform 1 0 18768 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_225
timestamp 1620791022
transform 1 0 21804 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_213
timestamp 1620791022
transform 1 0 20700 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_237
timestamp 1620791022
transform 1 0 22908 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_249
timestamp 1620791022
transform 1 0 24012 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_270
timestamp 1620791022
transform 1 0 25944 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_258
timestamp 1620791022
transform 1 0 24840 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1620791022
transform 1 0 24748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_282
timestamp 1620791022
transform 1 0 27048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_298
timestamp 1620791022
transform 1 0 28520 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_294
timestamp 1620791022
transform 1 0 28152 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1620791022
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1620791022
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1620791022
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1620791022
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1620791022
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1620791022
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_51
timestamp 1620791022
transform 1 0 5796 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_58
timestamp 1620791022
transform 1 0 6440 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1620791022
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_82
timestamp 1620791022
transform 1 0 8648 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_70
timestamp 1620791022
transform 1 0 7544 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_94
timestamp 1620791022
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1620791022
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1620791022
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_106
timestamp 1620791022
transform 1 0 10856 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_139
timestamp 1620791022
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_127
timestamp 1620791022
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_151
timestamp 1620791022
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_163
timestamp 1620791022
transform 1 0 16100 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1620791022
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1620791022
transform 1 0 16928 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1620791022
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1620791022
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1620791022
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1620791022
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1620791022
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_220
timestamp 1620791022
transform 1 0 21344 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_241
timestamp 1620791022
transform 1 0 23276 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_265
timestamp 1620791022
transform 1 0 25484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_253
timestamp 1620791022
transform 1 0 24380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_286
timestamp 1620791022
transform 1 0 27416 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1620791022
transform 1 0 27324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_277
timestamp 1620791022
transform 1 0 26588 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_298
timestamp 1620791022
transform 1 0 28520 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1620791022
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1620791022
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1620791022
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1620791022
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1620791022
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_30
timestamp 1620791022
transform 1 0 3864 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1620791022
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_54
timestamp 1620791022
transform 1 0 6072 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_42
timestamp 1620791022
transform 1 0 4968 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_66
timestamp 1620791022
transform 1 0 7176 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_78
timestamp 1620791022
transform 1 0 8280 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_99
timestamp 1620791022
transform 1 0 10212 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1620791022
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1620791022
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1620791022
transform 1 0 12420 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_111
timestamp 1620791022
transform 1 0 11316 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_144
timestamp 1620791022
transform 1 0 14352 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1620791022
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_135
timestamp 1620791022
transform 1 0 13524 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1620791022
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_180
timestamp 1620791022
transform 1 0 17664 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1620791022
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_201
timestamp 1620791022
transform 1 0 19596 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1620791022
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_192
timestamp 1620791022
transform 1 0 18768 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_225
timestamp 1620791022
transform 1 0 21804 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_213
timestamp 1620791022
transform 1 0 20700 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_237
timestamp 1620791022
transform 1 0 22908 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_249
timestamp 1620791022
transform 1 0 24012 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_270
timestamp 1620791022
transform 1 0 25944 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_258
timestamp 1620791022
transform 1 0 24840 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1620791022
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_282
timestamp 1620791022
transform 1 0 27048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_298
timestamp 1620791022
transform 1 0 28520 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_294
timestamp 1620791022
transform 1 0 28152 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1620791022
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1620791022
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1620791022
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1620791022
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1620791022
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1620791022
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1620791022
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1620791022
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_30
timestamp 1620791022
transform 1 0 3864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1620791022
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1620791022
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1620791022
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_51
timestamp 1620791022
transform 1 0 5796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_54
timestamp 1620791022
transform 1 0 6072 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_42
timestamp 1620791022
transform 1 0 4968 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_58
timestamp 1620791022
transform 1 0 6440 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1620791022
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1620791022
transform 1 0 7176 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_82
timestamp 1620791022
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_70
timestamp 1620791022
transform 1 0 7544 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_78
timestamp 1620791022
transform 1 0 8280 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_99
timestamp 1620791022
transform 1 0 10212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_87
timestamp 1620791022
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1620791022
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1620791022
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1620791022
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_111
timestamp 1620791022
transform 1 0 11316 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_115
timestamp 1620791022
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1620791022
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_106
timestamp 1620791022
transform 1 0 10856 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_144
timestamp 1620791022
transform 1 0 14352 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1620791022
transform 1 0 13892 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1620791022
transform 1 0 12788 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1620791022
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_135
timestamp 1620791022
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_156
timestamp 1620791022
transform 1 0 15456 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_151
timestamp 1620791022
transform 1 0 14996 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_163
timestamp 1620791022
transform 1 0 16100 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_180
timestamp 1620791022
transform 1 0 17664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_168
timestamp 1620791022
transform 1 0 16560 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1620791022
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1620791022
transform 1 0 16928 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1620791022
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1620791022
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1620791022
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1620791022
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1620791022
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_192
timestamp 1620791022
transform 1 0 18768 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_225
timestamp 1620791022
transform 1 0 21804 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_213
timestamp 1620791022
transform 1 0 20700 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_229
timestamp 1620791022
transform 1 0 22172 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1620791022
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_220
timestamp 1620791022
transform 1 0 21344 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_237
timestamp 1620791022
transform 1 0 22908 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_241
timestamp 1620791022
transform 1 0 23276 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_249
timestamp 1620791022
transform 1 0 24012 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_270
timestamp 1620791022
transform 1 0 25944 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_258
timestamp 1620791022
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_265
timestamp 1620791022
transform 1 0 25484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_253
timestamp 1620791022
transform 1 0 24380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1620791022
transform 1 0 24748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_282
timestamp 1620791022
transform 1 0 27048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_286
timestamp 1620791022
transform 1 0 27416 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1620791022
transform 1 0 27324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_277
timestamp 1620791022
transform 1 0 26588 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_298
timestamp 1620791022
transform 1 0 28520 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_298
timestamp 1620791022
transform 1 0 28520 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_294
timestamp 1620791022
transform 1 0 28152 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1620791022
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1620791022
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1620791022
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1620791022
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1620791022
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1620791022
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1620791022
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_51
timestamp 1620791022
transform 1 0 5796 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_58
timestamp 1620791022
transform 1 0 6440 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1620791022
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_82
timestamp 1620791022
transform 1 0 8648 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_70
timestamp 1620791022
transform 1 0 7544 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1620791022
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_115
timestamp 1620791022
transform 1 0 11684 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1620791022
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_106
timestamp 1620791022
transform 1 0 10856 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_139
timestamp 1620791022
transform 1 0 13892 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_127
timestamp 1620791022
transform 1 0 12788 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_151
timestamp 1620791022
transform 1 0 14996 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_163
timestamp 1620791022
transform 1 0 16100 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1620791022
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_172
timestamp 1620791022
transform 1 0 16928 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1620791022
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1620791022
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1620791022
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_229
timestamp 1620791022
transform 1 0 22172 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1620791022
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_220
timestamp 1620791022
transform 1 0 21344 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_241
timestamp 1620791022
transform 1 0 23276 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_265
timestamp 1620791022
transform 1 0 25484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_253
timestamp 1620791022
transform 1 0 24380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_286
timestamp 1620791022
transform 1 0 27416 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1620791022
transform 1 0 27324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_277
timestamp 1620791022
transform 1 0 26588 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1620791022
transform 1 0 28520 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1620791022
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1620791022
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1620791022
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1620791022
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1620791022
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_30
timestamp 1620791022
transform 1 0 3864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1620791022
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_54
timestamp 1620791022
transform 1 0 6072 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_42
timestamp 1620791022
transform 1 0 4968 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_66
timestamp 1620791022
transform 1 0 7176 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_78
timestamp 1620791022
transform 1 0 8280 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_99
timestamp 1620791022
transform 1 0 10212 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_87
timestamp 1620791022
transform 1 0 9108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1620791022
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_123
timestamp 1620791022
transform 1 0 12420 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_111
timestamp 1620791022
transform 1 0 11316 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_144
timestamp 1620791022
transform 1 0 14352 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1620791022
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_135
timestamp 1620791022
transform 1 0 13524 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1620791022
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_180
timestamp 1620791022
transform 1 0 17664 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1620791022
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1620791022
transform 1 0 19596 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1620791022
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_192
timestamp 1620791022
transform 1 0 18768 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_225
timestamp 1620791022
transform 1 0 21804 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_213
timestamp 1620791022
transform 1 0 20700 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_237
timestamp 1620791022
transform 1 0 22908 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_249
timestamp 1620791022
transform 1 0 24012 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_270
timestamp 1620791022
transform 1 0 25944 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1620791022
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1620791022
transform 1 0 24748 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_282
timestamp 1620791022
transform 1 0 27048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_298
timestamp 1620791022
transform 1 0 28520 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_294
timestamp 1620791022
transform 1 0 28152 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1620791022
transform -1 0 28888 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1620791022
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1620791022
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1620791022
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1620791022
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1620791022
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_51
timestamp 1620791022
transform 1 0 5796 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_58
timestamp 1620791022
transform 1 0 6440 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1620791022
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_82
timestamp 1620791022
transform 1 0 8648 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_70
timestamp 1620791022
transform 1 0 7544 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_94
timestamp 1620791022
transform 1 0 9752 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_115
timestamp 1620791022
transform 1 0 11684 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1620791022
transform 1 0 11592 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_106
timestamp 1620791022
transform 1 0 10856 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_139
timestamp 1620791022
transform 1 0 13892 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_127
timestamp 1620791022
transform 1 0 12788 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1620791022
transform 1 0 14996 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_163
timestamp 1620791022
transform 1 0 16100 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1620791022
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_172
timestamp 1620791022
transform 1 0 16928 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1620791022
transform 1 0 16836 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1620791022
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1620791022
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_229
timestamp 1620791022
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1620791022
transform 1 0 22080 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_220
timestamp 1620791022
transform 1 0 21344 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_241
timestamp 1620791022
transform 1 0 23276 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_265
timestamp 1620791022
transform 1 0 25484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_253
timestamp 1620791022
transform 1 0 24380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_286
timestamp 1620791022
transform 1 0 27416 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1620791022
transform 1 0 27324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_277
timestamp 1620791022
transform 1 0 26588 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_298
timestamp 1620791022
transform 1 0 28520 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1620791022
transform -1 0 28888 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1620791022
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1620791022
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1620791022
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1620791022
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_30
timestamp 1620791022
transform 1 0 3864 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1620791022
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_54
timestamp 1620791022
transform 1 0 6072 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_42
timestamp 1620791022
transform 1 0 4968 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_66
timestamp 1620791022
transform 1 0 7176 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_78
timestamp 1620791022
transform 1 0 8280 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_99
timestamp 1620791022
transform 1 0 10212 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_87
timestamp 1620791022
transform 1 0 9108 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1620791022
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_123
timestamp 1620791022
transform 1 0 12420 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_111
timestamp 1620791022
transform 1 0 11316 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_144
timestamp 1620791022
transform 1 0 14352 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1620791022
transform 1 0 14260 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_135
timestamp 1620791022
transform 1 0 13524 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_156
timestamp 1620791022
transform 1 0 15456 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_180
timestamp 1620791022
transform 1 0 17664 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_168
timestamp 1620791022
transform 1 0 16560 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_201
timestamp 1620791022
transform 1 0 19596 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1620791022
transform 1 0 19504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_192
timestamp 1620791022
transform 1 0 18768 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_225
timestamp 1620791022
transform 1 0 21804 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_213
timestamp 1620791022
transform 1 0 20700 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_237
timestamp 1620791022
transform 1 0 22908 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_249
timestamp 1620791022
transform 1 0 24012 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_270
timestamp 1620791022
transform 1 0 25944 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_258
timestamp 1620791022
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1620791022
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_282
timestamp 1620791022
transform 1 0 27048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_298
timestamp 1620791022
transform 1 0 28520 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_294
timestamp 1620791022
transform 1 0 28152 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1620791022
transform -1 0 28888 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1620791022
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1620791022
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1620791022
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1620791022
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1620791022
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1620791022
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_27
timestamp 1620791022
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_30
timestamp 1620791022
transform 1 0 3864 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1620791022
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1620791022
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1620791022
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_51
timestamp 1620791022
transform 1 0 5796 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_54
timestamp 1620791022
transform 1 0 6072 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_42
timestamp 1620791022
transform 1 0 4968 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_58
timestamp 1620791022
transform 1 0 6440 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1620791022
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_66
timestamp 1620791022
transform 1 0 7176 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_82
timestamp 1620791022
transform 1 0 8648 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_70
timestamp 1620791022
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_78
timestamp 1620791022
transform 1 0 8280 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_99
timestamp 1620791022
transform 1 0 10212 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_87
timestamp 1620791022
transform 1 0 9108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_94
timestamp 1620791022
transform 1 0 9752 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1620791022
transform 1 0 9016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_123
timestamp 1620791022
transform 1 0 12420 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_111
timestamp 1620791022
transform 1 0 11316 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_115
timestamp 1620791022
transform 1 0 11684 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1620791022
transform 1 0 11592 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_106
timestamp 1620791022
transform 1 0 10856 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_144
timestamp 1620791022
transform 1 0 14352 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_139
timestamp 1620791022
transform 1 0 13892 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_127
timestamp 1620791022
transform 1 0 12788 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1620791022
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_135
timestamp 1620791022
transform 1 0 13524 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_156
timestamp 1620791022
transform 1 0 15456 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_151
timestamp 1620791022
transform 1 0 14996 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_163
timestamp 1620791022
transform 1 0 16100 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_180
timestamp 1620791022
transform 1 0 17664 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_168
timestamp 1620791022
transform 1 0 16560 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1620791022
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_172
timestamp 1620791022
transform 1 0 16928 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1620791022
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_201
timestamp 1620791022
transform 1 0 19596 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1620791022
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1620791022
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1620791022
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_192
timestamp 1620791022
transform 1 0 18768 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_225
timestamp 1620791022
transform 1 0 21804 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_213
timestamp 1620791022
transform 1 0 20700 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_229
timestamp 1620791022
transform 1 0 22172 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1620791022
transform 1 0 22080 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_220
timestamp 1620791022
transform 1 0 21344 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_237
timestamp 1620791022
transform 1 0 22908 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_241
timestamp 1620791022
transform 1 0 23276 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_249
timestamp 1620791022
transform 1 0 24012 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_270
timestamp 1620791022
transform 1 0 25944 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_258
timestamp 1620791022
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_265
timestamp 1620791022
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_253
timestamp 1620791022
transform 1 0 24380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1620791022
transform 1 0 24748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_282
timestamp 1620791022
transform 1 0 27048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_286
timestamp 1620791022
transform 1 0 27416 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1620791022
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_277
timestamp 1620791022
transform 1 0 26588 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_298
timestamp 1620791022
transform 1 0 28520 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_298
timestamp 1620791022
transform 1 0 28520 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1620791022
transform 1 0 28152 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1620791022
transform -1 0 28888 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1620791022
transform -1 0 28888 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1620791022
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1620791022
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1620791022
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1620791022
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1620791022
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_51
timestamp 1620791022
transform 1 0 5796 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_58
timestamp 1620791022
transform 1 0 6440 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1620791022
transform 1 0 6348 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_82
timestamp 1620791022
transform 1 0 8648 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_70
timestamp 1620791022
transform 1 0 7544 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_94
timestamp 1620791022
transform 1 0 9752 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_115
timestamp 1620791022
transform 1 0 11684 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1620791022
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_106
timestamp 1620791022
transform 1 0 10856 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_139
timestamp 1620791022
transform 1 0 13892 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_127
timestamp 1620791022
transform 1 0 12788 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_151
timestamp 1620791022
transform 1 0 14996 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_163
timestamp 1620791022
transform 1 0 16100 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1620791022
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_172
timestamp 1620791022
transform 1 0 16928 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1620791022
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1620791022
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1620791022
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_229
timestamp 1620791022
transform 1 0 22172 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1620791022
transform 1 0 22080 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_220
timestamp 1620791022
transform 1 0 21344 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_241
timestamp 1620791022
transform 1 0 23276 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_265
timestamp 1620791022
transform 1 0 25484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_253
timestamp 1620791022
transform 1 0 24380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_286
timestamp 1620791022
transform 1 0 27416 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1620791022
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_277
timestamp 1620791022
transform 1 0 26588 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_298
timestamp 1620791022
transform 1 0 28520 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1620791022
transform -1 0 28888 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1620791022
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1620791022
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1620791022
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_27
timestamp 1620791022
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_30
timestamp 1620791022
transform 1 0 3864 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1620791022
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_54
timestamp 1620791022
transform 1 0 6072 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_42
timestamp 1620791022
transform 1 0 4968 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_66
timestamp 1620791022
transform 1 0 7176 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_78
timestamp 1620791022
transform 1 0 8280 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_99
timestamp 1620791022
transform 1 0 10212 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_87
timestamp 1620791022
transform 1 0 9108 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1620791022
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_123
timestamp 1620791022
transform 1 0 12420 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_111
timestamp 1620791022
transform 1 0 11316 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_144
timestamp 1620791022
transform 1 0 14352 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1620791022
transform 1 0 14260 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_135
timestamp 1620791022
transform 1 0 13524 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1620791022
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_180
timestamp 1620791022
transform 1 0 17664 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1620791022
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_201
timestamp 1620791022
transform 1 0 19596 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1620791022
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_192
timestamp 1620791022
transform 1 0 18768 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_225
timestamp 1620791022
transform 1 0 21804 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_213
timestamp 1620791022
transform 1 0 20700 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_237
timestamp 1620791022
transform 1 0 22908 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_249
timestamp 1620791022
transform 1 0 24012 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_270
timestamp 1620791022
transform 1 0 25944 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_258
timestamp 1620791022
transform 1 0 24840 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1620791022
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_282
timestamp 1620791022
transform 1 0 27048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_298
timestamp 1620791022
transform 1 0 28520 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_294
timestamp 1620791022
transform 1 0 28152 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1620791022
transform -1 0 28888 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1620791022
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1620791022
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1620791022
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1620791022
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1620791022
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_51
timestamp 1620791022
transform 1 0 5796 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_58
timestamp 1620791022
transform 1 0 6440 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1620791022
transform 1 0 6348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_82
timestamp 1620791022
transform 1 0 8648 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_70
timestamp 1620791022
transform 1 0 7544 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_94
timestamp 1620791022
transform 1 0 9752 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_115
timestamp 1620791022
transform 1 0 11684 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1620791022
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_106
timestamp 1620791022
transform 1 0 10856 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_139
timestamp 1620791022
transform 1 0 13892 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_127
timestamp 1620791022
transform 1 0 12788 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_151
timestamp 1620791022
transform 1 0 14996 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_163
timestamp 1620791022
transform 1 0 16100 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1620791022
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_172
timestamp 1620791022
transform 1 0 16928 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1620791022
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1620791022
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1620791022
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_229
timestamp 1620791022
transform 1 0 22172 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1620791022
transform 1 0 22080 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_220
timestamp 1620791022
transform 1 0 21344 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_241
timestamp 1620791022
transform 1 0 23276 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_265
timestamp 1620791022
transform 1 0 25484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_253
timestamp 1620791022
transform 1 0 24380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_286
timestamp 1620791022
transform 1 0 27416 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1620791022
transform 1 0 27324 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_277
timestamp 1620791022
transform 1 0 26588 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_298
timestamp 1620791022
transform 1 0 28520 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1620791022
transform -1 0 28888 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1620791022
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1620791022
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1620791022
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_27
timestamp 1620791022
transform 1 0 3588 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_30
timestamp 1620791022
transform 1 0 3864 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1620791022
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_54
timestamp 1620791022
transform 1 0 6072 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_42
timestamp 1620791022
transform 1 0 4968 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_66
timestamp 1620791022
transform 1 0 7176 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_78
timestamp 1620791022
transform 1 0 8280 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_99
timestamp 1620791022
transform 1 0 10212 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_87
timestamp 1620791022
transform 1 0 9108 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1620791022
transform 1 0 9016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_123
timestamp 1620791022
transform 1 0 12420 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_111
timestamp 1620791022
transform 1 0 11316 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_144
timestamp 1620791022
transform 1 0 14352 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1620791022
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_135
timestamp 1620791022
transform 1 0 13524 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_156
timestamp 1620791022
transform 1 0 15456 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_180
timestamp 1620791022
transform 1 0 17664 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_168
timestamp 1620791022
transform 1 0 16560 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_201
timestamp 1620791022
transform 1 0 19596 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1620791022
transform 1 0 19504 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_192
timestamp 1620791022
transform 1 0 18768 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_225
timestamp 1620791022
transform 1 0 21804 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_213
timestamp 1620791022
transform 1 0 20700 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_237
timestamp 1620791022
transform 1 0 22908 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_249
timestamp 1620791022
transform 1 0 24012 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_270
timestamp 1620791022
transform 1 0 25944 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_258
timestamp 1620791022
transform 1 0 24840 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1620791022
transform 1 0 24748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_282
timestamp 1620791022
transform 1 0 27048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_298
timestamp 1620791022
transform 1 0 28520 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_294
timestamp 1620791022
transform 1 0 28152 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1620791022
transform -1 0 28888 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1620791022
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1620791022
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1620791022
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1620791022
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1620791022
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_51
timestamp 1620791022
transform 1 0 5796 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_58
timestamp 1620791022
transform 1 0 6440 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1620791022
transform 1 0 6348 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_82
timestamp 1620791022
transform 1 0 8648 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_70
timestamp 1620791022
transform 1 0 7544 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_94
timestamp 1620791022
transform 1 0 9752 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_115
timestamp 1620791022
transform 1 0 11684 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1620791022
transform 1 0 11592 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_106
timestamp 1620791022
transform 1 0 10856 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_139
timestamp 1620791022
transform 1 0 13892 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_127
timestamp 1620791022
transform 1 0 12788 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_151
timestamp 1620791022
transform 1 0 14996 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_163
timestamp 1620791022
transform 1 0 16100 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1620791022
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_172
timestamp 1620791022
transform 1 0 16928 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1620791022
transform 1 0 16836 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1620791022
transform 1 0 20240 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1620791022
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_229
timestamp 1620791022
transform 1 0 22172 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1620791022
transform 1 0 22080 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_220
timestamp 1620791022
transform 1 0 21344 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_241
timestamp 1620791022
transform 1 0 23276 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_265
timestamp 1620791022
transform 1 0 25484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_253
timestamp 1620791022
transform 1 0 24380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_286
timestamp 1620791022
transform 1 0 27416 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1620791022
transform 1 0 27324 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_277
timestamp 1620791022
transform 1 0 26588 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_298
timestamp 1620791022
transform 1 0 28520 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1620791022
transform -1 0 28888 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1620791022
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1620791022
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1620791022
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1620791022
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1620791022
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1620791022
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_27
timestamp 1620791022
transform 1 0 3588 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1620791022
transform 1 0 4692 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1620791022
transform 1 0 3588 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_30
timestamp 1620791022
transform 1 0 3864 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1620791022
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_51
timestamp 1620791022
transform 1 0 5796 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_58
timestamp 1620791022
transform 1 0 6440 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_54
timestamp 1620791022
transform 1 0 6072 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_42
timestamp 1620791022
transform 1 0 4968 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1620791022
transform 1 0 6348 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_82
timestamp 1620791022
transform 1 0 8648 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_70
timestamp 1620791022
transform 1 0 7544 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_66
timestamp 1620791022
transform 1 0 7176 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_78
timestamp 1620791022
transform 1 0 8280 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_94
timestamp 1620791022
transform 1 0 9752 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_99
timestamp 1620791022
transform 1 0 10212 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_87
timestamp 1620791022
transform 1 0 9108 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1620791022
transform 1 0 9016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_115
timestamp 1620791022
transform 1 0 11684 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_123
timestamp 1620791022
transform 1 0 12420 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_111
timestamp 1620791022
transform 1 0 11316 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1620791022
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_106
timestamp 1620791022
transform 1 0 10856 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_139
timestamp 1620791022
transform 1 0 13892 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_127
timestamp 1620791022
transform 1 0 12788 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_144
timestamp 1620791022
transform 1 0 14352 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1620791022
transform 1 0 14260 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_135
timestamp 1620791022
transform 1 0 13524 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_151
timestamp 1620791022
transform 1 0 14996 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_156
timestamp 1620791022
transform 1 0 15456 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_163
timestamp 1620791022
transform 1 0 16100 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1620791022
transform 1 0 18032 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_172
timestamp 1620791022
transform 1 0 16928 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_180
timestamp 1620791022
transform 1 0 17664 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_168
timestamp 1620791022
transform 1 0 16560 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1620791022
transform 1 0 16836 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_208
timestamp 1620791022
transform 1 0 20240 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_196
timestamp 1620791022
transform 1 0 19136 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_201
timestamp 1620791022
transform 1 0 19596 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1620791022
transform 1 0 19504 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_192
timestamp 1620791022
transform 1 0 18768 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_229
timestamp 1620791022
transform 1 0 22172 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_225
timestamp 1620791022
transform 1 0 21804 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_213
timestamp 1620791022
transform 1 0 20700 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1620791022
transform 1 0 22080 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_220
timestamp 1620791022
transform 1 0 21344 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_241
timestamp 1620791022
transform 1 0 23276 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1620791022
transform 1 0 22908 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_249
timestamp 1620791022
transform 1 0 24012 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_265
timestamp 1620791022
transform 1 0 25484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_253
timestamp 1620791022
transform 1 0 24380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_270
timestamp 1620791022
transform 1 0 25944 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_258
timestamp 1620791022
transform 1 0 24840 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1620791022
transform 1 0 24748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_286
timestamp 1620791022
transform 1 0 27416 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_282
timestamp 1620791022
transform 1 0 27048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1620791022
transform 1 0 27324 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_277
timestamp 1620791022
transform 1 0 26588 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_298
timestamp 1620791022
transform 1 0 28520 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_298
timestamp 1620791022
transform 1 0 28520 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_294
timestamp 1620791022
transform 1 0 28152 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1620791022
transform -1 0 28888 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1620791022
transform -1 0 28888 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1620791022
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1620791022
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1620791022
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_27
timestamp 1620791022
transform 1 0 3588 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_30
timestamp 1620791022
transform 1 0 3864 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1620791022
transform 1 0 3772 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_54
timestamp 1620791022
transform 1 0 6072 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_42
timestamp 1620791022
transform 1 0 4968 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_66
timestamp 1620791022
transform 1 0 7176 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_78
timestamp 1620791022
transform 1 0 8280 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_99
timestamp 1620791022
transform 1 0 10212 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_87
timestamp 1620791022
transform 1 0 9108 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1620791022
transform 1 0 9016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_123
timestamp 1620791022
transform 1 0 12420 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_111
timestamp 1620791022
transform 1 0 11316 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_144
timestamp 1620791022
transform 1 0 14352 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1620791022
transform 1 0 14260 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_135
timestamp 1620791022
transform 1 0 13524 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_156
timestamp 1620791022
transform 1 0 15456 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_180
timestamp 1620791022
transform 1 0 17664 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_168
timestamp 1620791022
transform 1 0 16560 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_201
timestamp 1620791022
transform 1 0 19596 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1620791022
transform 1 0 19504 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_192
timestamp 1620791022
transform 1 0 18768 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_225
timestamp 1620791022
transform 1 0 21804 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_213
timestamp 1620791022
transform 1 0 20700 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_237
timestamp 1620791022
transform 1 0 22908 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_249
timestamp 1620791022
transform 1 0 24012 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_270
timestamp 1620791022
transform 1 0 25944 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_258
timestamp 1620791022
transform 1 0 24840 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1620791022
transform 1 0 24748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_282
timestamp 1620791022
transform 1 0 27048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_298
timestamp 1620791022
transform 1 0 28520 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_294
timestamp 1620791022
transform 1 0 28152 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1620791022
transform -1 0 28888 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1620791022
transform 1 0 2484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1620791022
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1620791022
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1620791022
transform 1 0 4692 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1620791022
transform 1 0 3588 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_51
timestamp 1620791022
transform 1 0 5796 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_58
timestamp 1620791022
transform 1 0 6440 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1620791022
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_82
timestamp 1620791022
transform 1 0 8648 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_70
timestamp 1620791022
transform 1 0 7544 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_94
timestamp 1620791022
transform 1 0 9752 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_115
timestamp 1620791022
transform 1 0 11684 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1620791022
transform 1 0 11592 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_106
timestamp 1620791022
transform 1 0 10856 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_139
timestamp 1620791022
transform 1 0 13892 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_127
timestamp 1620791022
transform 1 0 12788 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_151
timestamp 1620791022
transform 1 0 14996 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_163
timestamp 1620791022
transform 1 0 16100 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1620791022
transform 1 0 18032 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_172
timestamp 1620791022
transform 1 0 16928 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1620791022
transform 1 0 16836 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_208
timestamp 1620791022
transform 1 0 20240 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_196
timestamp 1620791022
transform 1 0 19136 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_229
timestamp 1620791022
transform 1 0 22172 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1620791022
transform 1 0 22080 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_220
timestamp 1620791022
transform 1 0 21344 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_241
timestamp 1620791022
transform 1 0 23276 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_265
timestamp 1620791022
transform 1 0 25484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_253
timestamp 1620791022
transform 1 0 24380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_286
timestamp 1620791022
transform 1 0 27416 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1620791022
transform 1 0 27324 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_277
timestamp 1620791022
transform 1 0 26588 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_298
timestamp 1620791022
transform 1 0 28520 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1620791022
transform -1 0 28888 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1620791022
transform 1 0 1380 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_6
timestamp 1620791022
transform 1 0 1656 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_18
timestamp 1620791022
transform 1 0 2760 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1620791022
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_30
timestamp 1620791022
transform 1 0 3864 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1620791022
transform 1 0 3772 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_26
timestamp 1620791022
transform 1 0 3496 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_59
timestamp 1620791022
transform 1 0 6532 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_42
timestamp 1620791022
transform 1 0 4968 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1620791022
transform 1 0 6440 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_54
timestamp 1620791022
transform 1 0 6072 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_71
timestamp 1620791022
transform 1 0 7636 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_83
timestamp 1620791022
transform 1 0 8740 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1620791022
transform 1 0 9568 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_95
timestamp 1620791022
transform 1 0 9844 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1620791022
transform 1 0 9108 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_88
timestamp 1620791022
transform 1 0 9200 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_115
timestamp 1620791022
transform 1 0 11684 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_117
timestamp 1620791022
transform 1 0 11868 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1620791022
transform 1 0 11776 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_107
timestamp 1620791022
transform 1 0 10948 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_129
timestamp 1620791022
transform 1 0 12972 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1620791022
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1620791022
transform 1 0 14076 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_158
timestamp 1620791022
transform 1 0 15640 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_146
timestamp 1620791022
transform 1 0 14536 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_175
timestamp 1620791022
transform 1 0 17204 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1620791022
transform 1 0 17112 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_170
timestamp 1620791022
transform 1 0 16744 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_187
timestamp 1620791022
transform 1 0 18308 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1620791022
transform -1 0 19412 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1620791022
transform 1 0 19044 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_204
timestamp 1620791022
transform 1 0 19872 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1620791022
transform 1 0 19780 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_199
timestamp 1620791022
transform 1 0 19412 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_216
timestamp 1620791022
transform 1 0 20976 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_228
timestamp 1620791022
transform 1 0 22080 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_245
timestamp 1620791022
transform 1 0 23644 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1620791022
transform 1 0 22540 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1620791022
transform 1 0 22448 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_262
timestamp 1620791022
transform 1 0 25208 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1620791022
transform 1 0 25116 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_257
timestamp 1620791022
transform 1 0 24748 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1620791022
transform 1 0 27784 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1620791022
transform -1 0 27416 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_286
timestamp 1620791022
transform 1 0 27416 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_291
timestamp 1620791022
transform 1 0 27876 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_274
timestamp 1620791022
transform 1 0 26312 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1620791022
transform -1 0 28888 0 -1 29920
box -38 -48 314 592
<< labels >>
rlabel metal2 s 10598 0 10654 800 6 clk
port 0 nsew signal input
rlabel metal2 s 19338 31368 19394 32168 6 l_sense
port 1 nsew signal input
rlabel metal2 s 9218 31368 9274 32168 6 l_thresh[0]
port 2 nsew signal input
rlabel metal2 s 478 0 534 800 6 l_thresh[1]
port 3 nsew signal input
rlabel metal2 s 29458 31368 29514 32168 6 m_sense
port 4 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 m_thresh_1
port 5 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 m_thresh_2
port 6 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 water_time_long
port 7 nsew signal input
rlabel metal3 s 29224 2048 30024 2168 6 water_time_short
port 8 nsew signal input
rlabel metal3 s 29224 17008 30024 17128 6 water_toggle
port 9 nsew signal tristate
rlabel metal4 s 24097 2128 24417 29968 6 VPWR
port 10 nsew power bidirectional
rlabel metal4 s 14836 2128 15156 29968 6 VPWR
port 11 nsew power bidirectional
rlabel metal4 s 5575 2128 5895 29968 6 VPWR
port 12 nsew power bidirectional
rlabel metal5 s 1104 25088 28888 25408 6 VPWR
port 13 nsew power bidirectional
rlabel metal5 s 1104 15840 28888 16160 6 VPWR
port 14 nsew power bidirectional
rlabel metal5 s 1104 6592 28888 6912 6 VPWR
port 15 nsew power bidirectional
rlabel metal4 s 19467 2128 19787 29968 6 VGND
port 16 nsew ground bidirectional
rlabel metal4 s 10205 2128 10525 29968 6 VGND
port 17 nsew ground bidirectional
rlabel metal5 s 1104 20464 28888 20784 6 VGND
port 18 nsew ground bidirectional
rlabel metal5 s 1104 11216 28888 11536 6 VGND
port 19 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30024 32168
<< end >>
