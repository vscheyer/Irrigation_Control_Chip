* SPICE3 file created from anADC.ext - technology: sky130A

.subckt sbc2 VP VN V1 V2 Vout nVout
X0 a_2280_320# a_3680_n450# nVout VN sky130_fd_pr__nfet_01v8 ad=1.5e+12p pd=8e+06u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X1 a_2060_n420# V1 a_760_n420# VN sky130_fd_pr__nfet_01v8 ad=1.5e+12p pd=8e+06u as=2.25e+12p ps=1.2e+07u w=1.5e+06u l=600000u
X2 a_1860_920# VP VP VP sky130_fd_pr__pfet_01v8 ad=3.75e+12p pd=2e+07u as=1.575e+13p ps=7.8e+07u w=1.5e+06u l=600000u
X3 a_320_320# a_100_n420# VP VP sky130_fd_pr__pfet_01v8 ad=3.75e+12p pd=2e+07u as=0p ps=0u w=1.5e+06u l=600000u
X4 VP VP a_100_320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X5 a_3680_n450# a_3680_n450# a_1860_920# VP sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=0p ps=0u w=1.5e+06u l=600000u
X6 VP VP a_1860_n1050# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X7 nVout a_3680_n450# a_2060_n420# VP sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X8 VP a_100_n420# a_2060_n420# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X9 VN a_100_320# a_320_n1050# VN sky130_fd_pr__nfet_01v8 ad=1.275e+13p pd=6.5e+07u as=3.75e+12p ps=2e+07u w=1.5e+06u l=600000u
X10 a_320_n1050# a_100_320# VP VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4.5e+12p ps=2.4e+07u w=1.5e+06u l=600000u
X11 a_320_n1050# a_100_320# VP VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X12 VN a_100_320# a_1860_n1050# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.75e+12p ps=2e+07u w=1.5e+06u l=600000u
X13 nVout a_3680_n450# a_2280_320# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X14 VN VN VP VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X15 a_320_320# a_100_n420# VN VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4.5e+12p ps=2.4e+07u w=1.5e+06u l=600000u
X16 VP a_100_n420# a_320_320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X17 a_100_n420# a_100_320# a_320_n1050# VN sky130_fd_pr__nfet_01v8 ad=1.5e+12p pd=8e+06u as=0p ps=0u w=1.5e+06u l=600000u
X18 Vout nVout VN VN sky130_fd_pr__nfet_01v8 ad=3e+12p pd=1.3e+07u as=0p ps=0u w=6e+06u l=150000u
X19 a_1860_n1050# a_3680_n450# a_3680_n450# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X20 a_1860_n1050# VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X21 a_2060_n420# VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X22 a_320_320# a_100_n420# VN VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X23 VP VP VN VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X24 Vout nVout VP VP sky130_fd_pr__pfet_01v8 ad=3e+12p pd=1.3e+07u as=0p ps=0u w=6e+06u l=150000u
X25 a_1860_920# VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X26 a_760_n420# a_100_320# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X27 a_320_n1050# a_100_320# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X28 VP a_100_320# a_320_n1050# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X29 a_100_320# a_100_n420# a_320_320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X30 a_2060_n420# a_3680_n450# nVout VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X31 VP a_100_320# a_320_n1050# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X32 a_1860_920# a_100_n420# a_100_n420# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X33 VP VP a_1860_920# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X34 VN VN a_100_n420# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X35 a_2060_n420# a_100_n420# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X36 a_100_320# VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X37 VN VN a_1860_n1050# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X38 VN a_100_n420# a_320_320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X39 VP VP a_1860_920# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X40 a_320_320# a_100_n420# a_100_320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X41 VN a_100_320# a_760_n420# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X42 a_1860_n1050# VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X43 a_320_n1050# a_100_320# VP VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X44 VP nVout Vout VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=150000u
X45 VN a_100_n420# a_320_320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X46 VN VN a_2060_n420# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X47 a_760_320# V1 a_2280_320# VP sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X48 a_1860_n1050# V2 a_2280_320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X49 VN VP VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X50 VP a_100_n420# a_1860_920# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X51 a_1860_920# a_3680_n450# a_3680_n450# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X52 a_3680_n450# a_3680_n450# a_1860_n1050# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X53 a_320_320# a_100_n420# VN VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X54 a_1860_920# a_100_n420# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X55 VP a_100_n420# a_760_320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X56 VN VN a_1860_n1050# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X57 a_2280_320# V2 a_1860_n1050# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X58 a_760_n420# V1 a_2060_n420# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X59 a_100_n420# a_100_n420# a_1860_920# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X60 a_2280_320# V1 a_760_320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X61 a_100_320# a_100_320# a_1860_n1050# VN sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=4e+06u as=0p ps=0u w=1.5e+06u l=600000u
X62 VN a_100_320# a_2280_320# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X63 a_760_n420# V2 a_1860_920# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X64 a_100_n420# VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X65 VN a_100_n420# a_320_320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X66 a_1860_920# V2 a_760_n420# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X67 VP a_100_320# a_320_n1050# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X68 a_1860_n1050# a_100_320# a_100_320# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X69 a_1860_n1050# a_100_320# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X70 a_760_320# a_100_n420# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X71 a_320_n1050# a_100_320# a_100_n420# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X72 VP VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X73 a_1860_n1050# VN VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X74 a_2280_320# a_100_320# VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
.ends

.subckt amux VP VN A B C Out
X0 VP C a_n50_680# VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X1 A C Out VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X2 Out C B VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X3 Out a_n50_680# B VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X4 A a_n50_680# Out VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X5 VN C a_n50_680# VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
.ends


* Top level circuit anADC

Xsbc2_0 VP VN sbc2_1/V1 OCC2 sbc2_0/Vout sbc2_0/nVout sbc2
Xsbc2_1 VP VN sbc2_1/V1 OCC1 OCC2 sbc2_1/nVout sbc2
Xsbc2_2 VP VN sbc2_2/V1 amux_1/A amux_1/A sbc2_2/nVout sbc2
Xamux_0 VP VN VL VH source amux_0/Out amux
Xamux_1 VP VN amux_1/A VN intc amux_1/Out amux
X0 a_n9470_n5530# a_1550_n5860# VN sky130_fd_pr__res_xhigh_po w=350000u l=5.29e+07u
X1 a_n8830_n4230# a_n4010_n4550# VN sky130_fd_pr__res_xhigh_po w=350000u l=2.19e+07u
X2 a_n8830_n3590# a_n4010_n3270# VN sky130_fd_pr__res_xhigh_po w=350000u l=2.19e+07u
X3 sbc2_1/V1 a_1550_n5200# VN sky130_fd_pr__res_xhigh_po w=350000u l=5.29e+07u
X4 Vtrip sbc2_0/Vout VN VN sky130_fd_pr__nfet_01v8 ad=1.5e+12p pd=7e+06u as=6.19e+12p ps=2.54e+07u w=3e+06u l=150000u
X5 sbc2_2/V1 a_n15480_n90# amux_0/Out VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X6 Vtrip sbc2_0/Vout VP VP sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=7e+06u as=2e+12p ps=1e+07u w=3e+06u l=150000u
X7 a_n20300_n5860# VN VN sky130_fd_pr__res_xhigh_po w=350000u l=4.85e+07u
X8 sbc2_2/V1 samp amux_0/Out VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X9 a_n8830_n2950# a_n4010_n2630# VN sky130_fd_pr__res_xhigh_po w=350000u l=2.19e+07u
X10 VP a_1550_n5860# VN sky130_fd_pr__res_xhigh_po w=350000u l=5.29e+07u
X11 sbc2_2/V1 VN sky130_fd_pr__cap_mim_m3_1 l=2e+07u w=2.5e+07u
X12 VP samp a_n15480_n90# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X13 OCC1 a_n4010_n2630# VN sky130_fd_pr__res_xhigh_po w=350000u l=2.19e+07u
X14 VN samp a_n15480_n90# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X15 amux_1/Out a_n4010_n4550# VN sky130_fd_pr__res_xhigh_po w=350000u l=2.19e+07u
X16 sbc2_1/nVout OCC2 sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2.5e+07u
X17 a_n8830_n3590# a_n4010_n3910# VN sky130_fd_pr__res_xhigh_po w=350000u l=2.19e+07u
X18 a_n20300_n5200# a_n10160_n5530# VN sky130_fd_pr__res_xhigh_po w=350000u l=4.85e+07u
X19 a_n20300_n5860# a_n10160_n5530# VN sky130_fd_pr__res_xhigh_po w=350000u l=4.85e+07u
X20 a_n20300_n5200# sbc2_1/V1 VN sky130_fd_pr__res_xhigh_po w=350000u l=4.85e+07u
X21 amux_1/A sbc2_2/nVout sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=2.5e+07u
X22 a_n8830_n4230# a_n4010_n3910# VN sky130_fd_pr__res_xhigh_po w=350000u l=2.19e+07u
X23 a_n8830_n2950# a_n4010_n3270# VN sky130_fd_pr__res_xhigh_po w=350000u l=2.19e+07u
X24 a_n9470_n5530# a_1550_n5200# VN sky130_fd_pr__res_xhigh_po w=350000u l=5.29e+07u
.end

